C0018801|033|heart failure
C0018801|033|hf
C0018801|033|congestive heart failure
C0018801|033|chf
C0018801|033|acute heart failure
C0018801|033|acute hf
C0018801|033|chronic heart failure
C0018801|033|chronic hf
C0018801|033|decompensated heart failure
C0018801|033|decompensated hf
C0018801|033|compensated heart failure
C0018801|033|compensated hf
C0018801|033|high-output heart failure
C0018801|033|low-output heart failure
C0018801|033|right heart failure
C0018801|033|right-sided heart failure
C0018801|033|right hf
C0018801|033|left heart failure
C0018801|033|left-sided heart failure
C0018801|033|left hf
C0018801|033|biventricular heart failure
C0018801|033|biventricular hf
C0018801|033|diastolic heart failure
C0018801|033|heart failure with preserved ejection fraction
C0018801|033|hfpef
C0018801|033|preserved ef heart failure
C0018801|033|systolic heart failure
C0018801|033|heart failure with reduced ejection fraction
C0018801|033|hfref
C0018801|033|reduced ef heart failure
C0018801|033|borderline ef heart failure
C0018801|033|mid-range ef heart failure
C0018801|033|hfmref
C0018801|033|ischemic heart failure
C0018801|033|ischemic hf
C0018801|033|nonischemic heart failure
C0018801|033|nonischemic hf
C0018801|033|valvular heart failure
C0018801|033|valvular hf
C0018801|033|hypertensive heart failure
C0018801|033|hypertensive hf
C0018801|033|amyloid heart failure
C0018801|033|amyloidosis-related hf
C0018801|033|cardiac amyloidosis with failure
C0018801|033|chemotherapy-induced heart failure
C0018801|033|chemo-induced hf
C0018801|033|peripartum cardiomyopathy
C0018801|033|tachycardia-induced heart failure
C0018801|033|tachycardia-induced hf
C0018801|033|myocarditis-induced heart failure
C0018801|033|myocarditis-related hf
C0018801|033|alcoholic cardiomyopathy with failure
C0018801|033|alcohol-related heart failure
C0018801|033|infiltrative cardiomyopathy with failure
C0018801|033|viral cardiomyopathy with failure
C0018801|033|postpartum heart failure
C0018801|033|dilated cardiomyopathy with failure
C0018801|033|dilated cm with hf
C0018801|033|idiopathic heart failure
C0018801|033|familial heart failure
C0018801|033|restrictive cardiomyopathy with failure
C0018801|033|rcm with hf
C0018801|033|cardiomyopathy with failure
C0018801|033|cm with hf
C0018801|033|advanced heart failure
C0018801|033|end-stage heart failure
C0018801|033|terminal heart failure
C0018801|033|refractory heart failure
C0018801|033|progressive heart failure
C0018801|033|acute on chronic heart failure
C0018801|033|aoc heart failure
C0018801|033|post-mi heart failure
C0018801|033|post-infarction heart failure
C0018801|033|cardiorenal syndrome
C0018801|033|pulmonary edema due to chf
C0018801|033|pump failure
C0018801|033|cardiac failure
C0018801|033|ventricular failure
C0018801|033|ventricular dysfunction
C0018801|033|lv failure
C0018801|033|left ventricular failure
C0018801|033|rv failure
C0018801|033|right ventricular failure
C0018801|033|congestive cardiac failure
C0018801|033|preload failure
C0018801|033|forward failure
C0018801|033|backward failure
C0018801|033|cardiac decompensation
C0018801|033|volume overload chf
C0018801|033|volume overload hf
C0018801|033|fluid overload chf
C0018801|033|fluid overload hf
C0018801|033|exacerbated chf
C0018801|033|exacerbation of hf
C0018801|033|cardiogenic pulmonary edema
C0018801|033|pulmonary congestion due to hf
C0018801|033|post-cardiac surgery hf
C0018801|033|iatrogenic heart failure
C0018801|033|drug-induced heart failure
C0018801|033|radiation-induced heart failure
C0018801|033|cor pulmonale with failure
C0018801|033|cor pulmonale with chf
C0018801|033|secondary heart failure
C0018801|033|primary heart failure
C0018801|033|tachyarrhythmia-related heart failure
C0018801|033|bradycardia-induced heart failure
C0018801|033|hfref exacerbation
C0018801|033|hfpef exacerbation
C0018801|033|heart failure with mid-range ef
C0018801|033|heart failure with mildly reduced ef
C0018801|033|diabetic cardiomyopathy with failure
C0018801|033|dm-related heart failure
C0018801|033|obesity-related heart failure
C0018801|033|thyrotoxic heart failure
C0018801|033|thyroid disease–related hf
C0018801|033|constrictive pericarditis with failure
C0018801|033|volume overloaded heart
C0018801|033|chf exacerbation
C0018801|033|new-onset heart failure
C0018801|033|new hf
C0018801|033|acute decompensated heart failure
C0018801|033|cardiac insufficiency
C0018801|033|chronic decompensated heart failure
C0018801|033|acute exacerbation of chf
C0018801|033|exertional heart failure
C0018801|033|post-viral heart failure
C0018801|033|post-viral cardiomyopathy with failure
C0018801|033|pericardial disease with failure
C0018801|033|transfusion-associated circulatory overload
C0018801|033|heart failure secondary to anemia
C0018801|033|high-output cardiac failure
C0018801|033|myocardial failure
C0018801|033|congestive myocardial failure
C0018801|033|acute left ventricular failure
C0018801|033|acute lvf
C0018801|033|chronic right heart failure
C0018801|033|heart failure with arrhythmia
C0018801|033|arrhythmia-related heart failure
C0018801|033|post-cardiotomy heart failure
C0018801|033|post-transplant heart failure
C0018801|033|transplant heart failure
C0018801|033|device-related heart failure
C0018801|033|lvad-related hf
C0018801|033|right heart dysfunction
C0018801|033|left heart dysfunction
C0018801|033|cardiac pump failure
C0018801|033|post-ischemic heart failure
C0018801|033|ischemic dilated cardiomyopathy with failure
C0018801|033|post-reperfusion heart failure
C0018801|033|stress-induced cardiomyopathy with failure
C0018801|033|takotsubo with failure
C0018801|033|takotsubo hf
C0018801|033|chagas disease with heart failure
C0018801|033|hereditary heart failure
C0018801|033|arvc with failure
C0018801|033|arrhythmogenic rv cardiomyopathy with hf
C0027051|033|myocardial infarction
C0027051|033|mi
C0027051|033|acute mi
C0027051|033|ami
C0027051|033|acute myocardial infarction
C0027051|033|stemi
C0027051|033|st-elevation mi
C0027051|033|st-elevation myocardial infarction
C0027051|033|nstemi
C0027051|033|non-st-elevation mi
C0027051|033|non-st-elevation myocardial infarction
C0027051|033|transmural mi
C0027051|033|subendocardial mi
C0027051|033|inferior mi
C0027051|033|anterior mi
C0027051|033|lateral mi
C0027051|033|posterior mi
C0027051|033|septal mi
C0027051|033|high lateral mi
C0027051|033|unstable coronary syndrome
C0027051|033|ischemic mi
C0027051|033|ischemic infarct
C0027051|033|cardiac infarct
C0027051|033|acute coronary syndrome
C0027051|033|acs
C0027051|033|coronary thrombosis
C0027051|033|coronary occlusion
C0027051|033|transmural infarct
C0027051|033|subendocardial infarct
C0027051|033|heart attack
C0027051|033|old mi
C0027051|033|prior mi
C0027051|033|healed mi
C0027051|033|silent infarction
C0027051|033|silent mi
C0027051|033|q wave mi
C0027051|033|non-q wave mi
C0027051|033|spontaneous mi
C0027051|033|type 1 mi
C0027051|033|type i mi
C0027051|033|type 2 mi
C0027051|033|type ii mi
C0027051|033|demand mi
C0027051|033|supply-demand mismatch mi
C0027051|033|secondary mi
C0027051|033|perioperative mi
C0027051|033|post-procedure mi
C0027051|033|stent thrombosis mi
C0027051|033|in-stent mi
C0027051|033|valvular mi
C0027051|033|hypertensive mi
C0027051|033|amyloid mi
C0027051|033|chemo-induced mi
C0027051|033|cancer therapy–related mi
C0027051|033|ppcm-related mi
C0027051|033|post-partum cm with mi
C0027051|033|myocarditis-related mi
C0027051|033|tachycardia-induced mi
C0027051|033|atrial fibrillation mi
C0027051|033|coronary embolism mi
C0027051|033|embolism-related mi
C0027051|033|coronary spasm mi
C0027051|033|vasospastic mi
C0027051|033|coronary dissection mi
C0027051|033|scad mi
C0027051|033|spontaneous coronary artery dissection mi
C0027051|033|thrombotic mi
C0027051|033|microvascular mi
C0027051|033|microvascular infarction
C0027051|033|cardiac necrosis
C0027051|033|myocardial necrosis
C0027051|033|myocardial injury (ischemic)
C0027051|033|ischemia-induced necrosis
C0027051|033|supply-demand mismatch infarct
C0027051|033|lv infarct
C0027051|033|rv infarct
C0027051|033|presumed mi
C0027051|033|possible mi
C0027051|033|probable mi
C0027051|033|unrecognized mi
C0027051|033|nontransmural mi
C0027051|033|recurrent mi
C0027051|033|multiple mi
C0027051|033|re-infarction
C0027051|033|reinfarction
C0027051|033|reinfarct
C0027051|033|reinfarcted myocardium
C0027051|033|extensive mi
C0027051|033|widespread mi
C0027051|033|limited mi
C0027051|033|microscopic mi
C0027051|033|multi-territory mi
C0027051|033|multivessel mi
C0027051|033|single vessel mi
C0027051|033|inferolateral mi
C0027051|033|anterolateral mi
C0027051|033|posterolateral mi
C0027051|033|apical mi
C0027051|033|basal mi
C0027051|033|old inferior mi
C0027051|033|old anterior mi
C0027051|033|old lateral mi
C0027051|033|old septal mi
C0027051|033|old transmural mi
C0027051|033|old subendocardial mi
C0027051|033|silent anterior mi
C0027051|033|silent inferior mi
C0027051|033|silent posterior mi
C0027051|033|acute infarct
C0027051|033|acute transmural mi
C0027051|033|acute subendocardial mi
C0027051|033|acute anterior mi
C0027051|033|acute inferior mi
C0027051|033|acute lateral mi
C0027051|033|acute septal mi
C0027051|033|acute posterior mi
C0027051|033|nstemi acs
C0027051|033|stemi acs
C0027051|033|post-cath mi
C0027051|033|periprocedural mi
C0027051|033|high sensitivity troponin mi
C0027051|033|troponin-positive mi
C0027051|033|troponin rise (mi)
C0027051|033|ihd with mi
C0027051|033|ischemic heart disease with mi
C0027051|033|cad with mi
C0027051|033|coronary artery disease with mi
C0027051|033|mi with lv dysfunction
C0027051|033|mi with heart failure
C0027051|033|chf secondary to mi
C0027051|033|ventricular infarct
C0027051|033|coronary syndrome (mi)
C0027051|033|infarcted myocardium
C0027051|033|myocardial infarct tissue
C0027051|033|fibrotic myocardium post mi
C0027051|033|scarred myocardium (post mi)
C0027051|033|cardiac event (infarct)
C0027051|033|myocardial event (inf. type)
C0027051|033|myocardial ischemia with infarction
C0027051|033|ischemic cardiomyopathy (mi)
C0027051|033|mi secondary to embolus
C0027051|033|mi secondary to spasm
C0027051|033|mi secondary to amyloid
C0027051|033|mi secondary to hypotension
C0027051|033|mi secondary to vasospasm
C0027051|033|mi secondary to thrombosis
C0027051|033|mi secondary to hypertension
C0027051|033|mi secondary to cocaine
C0027051|033|cocaine-induced mi
C0027051|033|mi secondary to anemia
C0027051|033|demand ischemia with infarct
C0027051|033|coronary supply mi
C0027051|033|coronary demand mi
C0027051|033|type 3 mi
C0027051|033|type iii mi
C0027051|033|type 4a mi
C0027051|033|type 4b mi
C0027051|033|type 4c mi
C0027051|033|type 5 mi
C0027051|033|post-pci mi
C0027051|033|post-cabg mi
C0027051|033|late mi
C0027051|033|early mi
C0027051|033|periinfarct
C0027051|033|myocardial infarct zone
C0027051|033|mi territory
C0027051|033|coronary syndrome (with mi)
C0027051|033|infarct-related artery
C0027051|033|culprit lesion mi
C0027051|033|mi with papillary muscle involvement
C0027051|033|acute infarction event
C0027051|033|cardiac event (mi type)
C0027051|033|coronary syndrome with infarct
C0027051|033|cardiac ischemic event
C0027051|033|acute plaque rupture mi
C0027051|033|mi with thrombus
C0002965|033|unstable angina
C0002965|033|ua
C0002965|033|acs-ua
C0002965|033|pre-infarction angina
C0002965|033|crescendo angina
C0002965|033|intermediate coronary syndrome
C0002965|033|preinfarction angina
C0002965|033|threatened mi
C0002965|033|angina at rest
C0002965|033|rest angina
C0002965|033|ischemic ua
C0002965|033|ischemic unstable angina
C0002965|033|acute isch angina
C0002965|033|non-st elevation acs-ua
C0002965|033|nstemi/ua
C0002965|033|nstemi rule out
C0002965|033|nstemi suspected/ua
C0002965|033|decubitus ua
C0002965|033|variant ua
C0002965|033|refractory ua
C0002965|033|angina exacerbation
C0002965|033|progressive angina
C0002965|033|worsening angina
C0002965|033|dynamic angina
C0002965|033|unstable exertional angina
C0002965|033|secondary unstable angina
C0002965|033|valvular ua
C0002965|033|valvular unstable angina
C0002965|033|hypertensive ua
C0002965|033|hypertensive unstable angina
C0002965|033|chemo-induced unstable angina
C0002965|033|drug-induced ua
C0002965|033|myocarditis-associated ua
C0002965|033|tachycardia-induced ua
C0002965|033|ppcm with ua
C0002965|033|nonischemic ua
C0002965|033|postintervention ua
C0002965|033|post-pci ua
C0002965|033|post-cabg ua
C0002965|033|bypass ua
C0002965|033|stent ua
C0002965|033|spontaneous unstable angina
C0002965|033|recurrent ua
C0002965|033|recurring unstable angina
C0002965|033|intractable ua
C0002965|033|resistant unstable angina
C0002965|033|unstable post-infarct angina
C0002965|033|angina instable
C0002965|033|instable angina
C0002965|033|angor instable
C0002965|033|ua/nstemi
C0002965|033|non-q-wave ua
C0002965|033|noq ua
C0002965|033|unstable ep angina
C0002965|033|ua w/elevated troponin
C0002965|033|ua (tn-)
C0038454|033|cerebrovascular accident
C0038454|033|cva
C0038454|033|stroke
C0038454|033|acute stroke
C0038454|033|embolic stroke
C0038454|033|thrombotic stroke
C0038454|033|hemorrhagic stroke
C0038454|033|ischemic stroke
C0038454|033|nonischemic stroke
C0038454|033|lacunar stroke
C0038454|033|cerebral infarct
C0038454|033|cerebral infarction
C0038454|033|cerebral hemorrhage
C0038454|033|brain attack
C0038454|033|brain infarct
C0038454|033|brain infarction
C0038454|033|acute cerebral infarct
C0038454|033|large vessel stroke
C0038454|033|small vessel stroke
C0038454|033|cryptogenic stroke
C0038454|033|watershed infarct
C0038454|033|tia with infarct
C0038454|033|intraparenchymal hemorrhage
C0038454|033|parenchymal hemorrhage
C0038454|033|icvh
C0038454|033|ich
C0038454|033|intracerebral hemorrhage
C0038454|033|subcortical infarct
C0038454|033|cortical infarct
C0038454|033|pca stroke
C0038454|033|mca stroke
C0038454|033|aca stroke
C0038454|033|posterior stroke
C0038454|033|anterior circulation stroke
C0038454|033|posterior circulation stroke
C0038454|033|valvular embolic stroke
C0038454|033|cardioembolic stroke
C0038454|033|atrial fib stroke
C0038454|033|afib stroke
C0038454|033|non-valvular stroke
C0038454|033|artery-to-artery embolic stroke
C0038454|033|arterial embolic stroke
C0038454|033|vertebrobasilar stroke
C0038454|033|basilar stroke
C0038454|033|brainstem stroke
C0038454|033|pontine stroke
C0038454|033|cerebellar stroke
C0038454|033|subarachnoid hemorrhage
C0038454|033|sah
C0038454|033|midline cerebral infarct
C0038454|033|right mca stroke
C0038454|033|left mca stroke
C0038454|033|r mca infarct
C0038454|033|l mca infarct
C0038454|033|left hemisphere infarct
C0038454|033|right hemisphere infarct
C0038454|033|r cortical stroke
C0038454|033|l cortical stroke
C0038454|033|chronic infarct
C0038454|033|acute on chronic infarct
C0038454|033|microvascular infarct
C0038454|033|silent infarct
C0038454|033|old infarct
C0038454|033|remote infarct
C0038454|033|multi-infarct
C0038454|033|multiple infarcts
C0038454|033|multi-territorial stroke
C0038454|033|transient cerebral ischemia
C0038454|033|cerebral ischemia
C0038454|033|acute cerebral ischemia
C0038454|033|territorial infarct
C0038454|033|territorial stroke
C0038454|033|territorial hemorrhage
C0038454|033|flow-related infarct
C0038454|033|global cerebral ischemia
C0038454|033|atherothrombotic stroke
C0038454|033|cholesterol embolic stroke
C0038454|033|calcific embolic stroke
C0038454|033|infective embolic stroke
C0038454|033|meningovascular stroke
C0038454|033|arteriopathic stroke
C0038454|033|hypertensive stroke
C0038454|033|hypertensive intracerebral hemorrhage
C0038454|033|amyloid angiopathy stroke
C0038454|033|amyloid angiopathy hemorrhage
C0038454|033|caa-associated hemorrhage
C0038454|033|leukoaraiosis-associated stroke
C0038454|033|chemo-induced stroke
C0038454|033|radiation-induced stroke
C0038454|033|drug-induced stroke
C0038454|033|ppcm-related stroke
C0038454|033|peripartum stroke
C0038454|033|pregnancy-associated stroke
C0038454|033|puerperal stroke
C0038454|033|myocarditis-associated stroke
C0038454|033|tachycardia-induced stroke
C0038454|033|arrhythmic embolic stroke
C0038454|033|endocarditis embolic stroke
C0038454|033|paradoxical embolic stroke
C0038454|033|nonbacterial thrombotic embolic stroke
C0038454|033|nbte stroke
C0038454|033|moya moya stroke
C0038454|033|vasculitis-associated stroke
C0038454|033|sle-associated stroke
C0038454|033|antiphospholipid stroke
C0038454|033|hypercoagulable stroke
C0038454|033|coagulopathy stroke
C0038454|033|cocaine-induced stroke
C0038454|033|vasospasm-associated infarct
C0038454|033|hypoperfusion stroke
C0038454|033|hemodynamic stroke
C0038454|033|low-flow infarct
C0038454|033|occlusive stroke
C0038454|033|arterial occlusive infarct
C0038454|033|arterial occlusion stroke
C0038454|033|large artery atherosclerotic stroke
C0038454|033|laa stroke
C0038454|033|intracranial atherosclerotic stroke
C0038454|033|extracranial atherosclerotic stroke
C0038454|033|atherothrombotic infarct
C0038454|033|cavitary infarct
C0038454|033|cavitating infarct
C0038454|033|encephalomalacic infarct
C0038454|033|encephalomalacia from cva
C0038454|033|cerebellar infarct
C0038454|033|cerebellar hemorrhage
C0038454|033|medullary infarct
C0038454|033|medullary stroke
C0038454|033|brainstem infarct
C0038454|033|thalamic infarct
C0038454|033|thalamic hemorrhage
C0038454|033|putaminal hemorrhage
C0038454|033|putaminal infarct
C0038454|033|capsular stroke
C0038454|033|internal capsule infarct
C0038454|033|subcortical hemorrhage
C0038454|033|subcortical stroke
C0038454|033|watershed stroke
C0038454|033|borderzone infarct
C0038454|033|lacunar infarct
C0038454|033|peri-ictal infarct
C0038454|033|hypoxic ischemic stroke
C0038454|033|cardiac arrest-related stroke
C0038454|033|post-cardiac arrest infarct
C0038454|033|cerebral embolism
C0038454|033|cerebral embolic event
C0038454|033|cerebral thromboembolism
C0038454|033|cerebrovascular event
C0038454|033|acute cerebrovascular event
C0038454|033|major stroke
C0038454|033|minor stroke
C0038454|033|silent stroke
C0038454|033|subclinical stroke
C0038454|033|cerebral event
C0038454|033|pres-associated infarct
C0038454|033|posterior reversible encephalopathy stroke
C0038454|033|arteriopathy-associated infarct
C0038454|033|cortical laminar necrosis
C0038454|033|subdural hematoma stroke
C0038454|033|cortical microinfarct
C0038454|033|cortical microbleed associated stroke
C0038454|033|embolism to brain
C0038454|033|embolus to brain
C0038454|033|cerebral occlusion event
C0038454|033|cerebral arterial infarct
C0038454|033|cerebral embologenic event
C0038454|033|left hemispheric stroke
C0038454|033|right hemispheric stroke
C0038454|033|left parietal stroke
C0038454|033|right parietal stroke
C0038454|033|left frontal infarct
C0038454|033|right frontal infarct
C0004238|033|atrial fibrillation
C0004238|033|af
C0004238|033|afib
C0004238|033|a-fib
C0004238|033|a fibrillation
C0004238|033|chronic atrial fibrillation
C0004238|033|paroxysmal atrial fibrillation
C0004238|033|persistent atrial fibrillation
C0004238|033|permanent atrial fibrillation
C0004238|033|long-standing persistent atrial fibrillation
C0004238|033|valvular atrial fibrillation
C0004238|033|nonvalvular atrial fibrillation
C0004238|033|nvaf
C0004238|033|valvular af
C0004238|033|nonvalvular af
C0004238|033|secondary atrial fibrillation
C0004238|033|recurrent atrial fibrillation
C0004238|033|acute atrial fibrillation
C0004238|033|postoperative atrial fibrillation
C0004238|033|new-onset atrial fibrillation
C0004238|033|lone atrial fibrillation
C0004238|033|ischemic atrial fibrillation
C0004238|033|nonischemic atrial fibrillation
C0004238|033|hypertensive atrial fibrillation
C0004238|033|amyloid atrial fibrillation
C0004238|033|amyloidosis-related af
C0004238|033|chemo-induced atrial fibrillation
C0004238|033|chemotherapy-related af
C0004238|033|tachycardia-induced atrial fibrillation
C0004238|033|tachy-induced af
C0004238|033|ppcm-related atrial fibrillation
C0004238|033|peripartum af
C0004238|033|myocarditis-associated af
C0004238|033|alcoholic af
C0004238|033|holiday heart syndrome
C0004238|033|alcohol-induced atrial fibrillation
C0004238|033|af with rvr
C0004238|033|atrial fibrillation with rapid ventricular response
C0004238|033|af w/ rvr
C0004238|033|af with slow ventricular response
C0004238|033|af with bradycardia
C0004238|033|subclinical atrial fibrillation
C0004238|033|asymptomatic atrial fibrillation
C0004238|033|symptomatic atrial fibrillation
C0004238|033|atrial fib
C0004238|033|atrial-fib
C0004238|033|fib/flutter
C0004238|033|af/flutter
C0004238|033|af/afl
C0004238|033|a fib/flutter
C0004238|033|paroxysmal af
C0004238|033|persistent af
C0004238|033|permanent af
C0004238|033|long-standing persistent af
C0004238|033|recurrent af
C0004238|033|secondary af
C0004238|033|acute af
C0004238|033|new-onset af
C0004238|033|postop af
C0004238|033|post-op af
C0004238|033|common-type atrial fibrillation
C0004238|033|rapid atrial fibrillation
C0004238|033|atrial fibrillation crisis
C0004238|033|resistant atrial fibrillation
C0004238|033|uncontrolled atrial fibrillation
C0004238|033|controlled atrial fibrillation
C0004238|033|a. fib.
C0004238|033|a/f
C0004238|033|a-fibrillation
C0004238|033|afib p/w rvr
C0004238|033|paroxysmal a-fib
C0004238|033|persistent a-fib
C0004238|033|permanent a-fib
C0004238|033|af with slow vr
C0004238|033|af w/ svr
C0004238|033|valvular a-fib
C0004238|033|nonvalvular a-fib
C0004238|033|non-ischemic af
C0004238|033|ischemic af
C0004238|033|hypertensive af
C0004238|033|ms/af
C0004238|033|mitral stenosis af
C0004238|033|rheumatic af
C0004238|033|chf with af
C0004238|033|hfpef with af
C0004238|033|hfref with af
C0004238|033|chf/af
C0004238|033|hf/af
C0004238|033|dilated cardiomyopathy with af
C0004238|033|dcm/af
C0004238|033|cardioembolic af
C0004238|033|thromboembolic af
C0004238|033|thyrotoxic af
C0004238|033|hyperthyroid af
C0004238|033|thyrotoxic atrial fibrillation
C0004238|033|post-cardiac surgery af
C0004238|033|surgery-induced af
C0004238|033|postablation af
C0004238|033|post-ablation a-fib
C0004238|033|lone af
C0004238|033|cryptogenic af
C0004238|033|familial af
C0004238|033|inherited af
C0004238|033|idiopathic af
C0004238|033|spontaneous af
C0004238|033|secondary to sepsis af
C0004238|033|sepsis-associated af
C0004238|033|post-mi af
C0004238|033|post infarct af
C0004238|033|post cabg af
C0004238|033|cabg-related af
C0004238|033|post-op a-fib
C0004238|033|perioperative af
C0004238|033|renal failure with af
C0004238|033|af in ckd
C0004238|033|esrd with af
C0004238|033|dialysis-associated af
C0004238|033|copd-related af
C0004238|033|obstructive sleep apnea with af
C0004238|033|osa with af
C0004238|033|af in elderly
C0004238|033|degenerative af
C0004238|033|afiv
C0004238|033|a fib
C0004238|033|afib episode
C0004238|033|asx af
C0004238|033|parox af
C0004238|033|sym af
C0004238|033|asymp af
C0004238|033|atrial fib episode
C0004238|033|beta-blocker controlled af
C0004238|033|rate-controlled af
C0004238|033|rhythm-controlled af
C0004238|033|af on anticoagulation
C0004238|033|af on oac
C0004238|033|af with stroke
C0004238|033|af with embolism
C0004238|033|embolic a-fib
C0004238|033|af of unknown cause
C0004238|033|af post anaesthesia
C0004238|033|af on ecg
C0004238|033|ecg: af
C0004238|033|telemetry: af
C0004238|033|holter: af
C0004238|033|atrial fib rvr
C0004238|033|fib w/ rvr
C0004238|033|af/svr
C0004238|033|tachy af
C0004238|033|persistent afib
C0004238|033|chronic afib
C0004238|033|recurring afib
C0004238|033|long-term afib
C0004238|033|persistent a fib
C0004238|033|intermittent af
C0004238|033|episodes of af
C0004238|033|brief af
C0004238|033|asx atrial fib
C0004238|033|supraventricular af
C0015672|033|fatigue
C0015672|033|fatigued
C0015672|033|fatiging
C0015672|033|fatigability
C0015672|033|easy fatigability
C0015672|033|early fatigability
C0015672|033|increased fatigability
C0015672|033|severe fatigue
C0015672|033|chronic fatigue
C0015672|033|malaise
C0015672|033|lassitude
C0015672|033|tired
C0015672|033|tiredness
C0015672|033|easily tired
C0015672|033|exercise intolerance
C0015672|033|dec exercise tolerance
C0015672|033|poor exercise tolerance
C0015672|033|exertional fatigue
C0015672|033|exercise-induced fatigue
C0015672|033|post-exertional fatigue
C0015672|033|weakness
C0015672|033|generalized weakness
C0015672|033|muscle weakness
C0015672|033|subjective weakness
C0015672|033|lethargy
C0015672|033|lethargic
C0015672|033|exhaustion
C0015672|033|exhausted
C0015672|033|low energy
C0015672|033|decreased energy
C0015672|033|dec energy
C0015672|033|loss of energy
C0015672|033|easy exhaustion
C0015672|033|quickly exhausted
C0015672|033|no stamina
C0015672|033|reduced stamina
C0015672|033|low stamina
C0015672|033|weariness
C0015672|033|worn out
C0015672|033|drained
C0015672|033|sluggishness
C0015672|033|sluggish
C0015672|033|slowness
C0015672|033|nonrestorative sleep
C0015672|033|non-restful sleep
C0015672|033|daytime sleepiness
C0015672|033|somnolence
C0015672|033|drowsiness
C0015672|033|sleepiness
C0015672|033|poor tolerance to activity
C0015672|033|activity intolerance
C0015672|033|easy fatigued
C0015672|033|subjective fatigue
C0015672|033|chemo-induced fatigue
C0015672|033|chemotherapy-related fatigue
C0015672|033|ca fatigue
C0015672|033|post-chemo fatigue
C0015672|033|cancer fatigue
C0015672|033|radiation-induced fatigue
C0015672|033|anemia-associated fatigue
C0015672|033|anemic fatigue
C0015672|033|hf fatigue
C0015672|033|chf fatigue
C0015672|033|heart failure fatigue
C0015672|033|ischemic fatigue
C0015672|033|low cardiac output fatigue
C0015672|033|amyloid fatigue
C0015672|033|amyloidosis-related fatigue
C0015672|033|valvular fatigue
C0015672|033|hypertensive fatigue
C0015672|033|htn fatigue
C0015672|033|htn-related fatigue
C0015672|033|myocarditis fatigue
C0015672|033|tachycardia-induced fatigue
C0015672|033|arrhythmia-related fatigue
C0015672|033|postviral fatigue
C0015672|033|viral fatigue
C0015672|033|infectious fatigue
C0015672|033|post-covid fatigue
C0015672|033|covid fatigue
C0015672|033|me/cfs
C0015672|033|chronic fatigue syndrome
C0015672|033|post-infectious fatigue
C0015672|033|hiv-related fatigue
C0015672|033|apls fatigue
C0015672|033|ppcm fatigue
C0015672|033|peripartum fatigue
C0015672|033|pregnancy-induced fatigue
C0015672|033|postpartum fatigue
C0015672|033|endocrine fatigue
C0015672|033|thyroid-related fatigue
C0015672|033|hypothyroid fatigue
C0015672|033|hypothyroidism fatigue
C0015672|033|adrenal fatigue
C0015672|033|addison’s fatigue
C0015672|033|diabetic fatigue
C0015672|033|renal fatigue
C0015672|033|ckd fatigue
C0015672|033|renal failure fatigue
C0015672|033|hepatic fatigue
C0015672|033|liver failure fatigue
C0015672|033|cld fatigue
C0015672|033|malignancy fatigue
C0015672|033|sle fatigue
C0015672|033|ra fatigue
C0015672|033|ms fatigue
C0015672|033|neuromuscular fatigue
C0015672|033|depression-related fatigue
C0015672|033|psychogenic fatigue
C0015672|033|mental fatigue
C0015672|033|cognitive fatigue
C0015672|033|fibromyalgia fatigue
C0015672|033|pain-related fatigue
C0015672|033|post-concussion fatigue
C0015672|033|tbi fatigue
C0015672|033|chronic disease fatigue
C0015672|033|post-surgical fatigue
C0015672|033|post-op fatigue
C0015672|033|drug-induced fatigue
C0015672|033|medication-related fatigue
C0015672|033|antidepressant fatigue
C0015672|033|antipsychotic fatigue
C0015672|033|sleep apnea fatigue
C0015672|033|osa fatigue
C0015672|033|csa fatigue
C0015672|033|night sweats and fatigue
C0015672|033|migrainous fatigue
C0015672|033|fatigue of unknown etiology
C0015672|033|idiopathic fatigue
C0015672|033|ebv fatigue
C0015672|033|lyme fatigue
C0015672|033|rheumatologic fatigue
C0015672|033|crps fatigue
C0015672|033|copd fatigue
C0015672|033|pulmonary fatigue
C0015672|033|respiratory fatigue
C0015672|033|disease-related fatigue
C0015672|033|tired out
C0015672|033|wiped out
C0015672|033|run down
C0015672|033|flagging
C0015672|033|lack of pep
C0015672|033|lack of vigor
C0015672|033|slowed down
C0015672|033|lacks energy
C0015672|033|needs naps
C0015672|033|falls asleep during day
C0015672|033|reduced activity tolerance
C0015672|033|reduced functional capacity
C0015672|033|cannot keep up usual activity
C0015672|033|mental exhaustion
C0015672|033|physical exhaustion
C0015672|033|overwhelming fatigue
C0015672|033|burnout
C0015672|033|asthenia
C0015672|033|listlessness
C0015672|033|debilitation
C0015672|033|debilitated
C0015672|033|profound fatigue
C0015672|033|significant fatigue
C0015672|033|marked fatigue
C0015672|033|extreme fatigue
C0015672|033|incapacitating fatigue
C0015672|033|insufficient energy
C0015672|033|difficulty completing tasks
C0015672|033|reports fatigue
C0015672|033|pt c/o fatigue
C0015672|033|c/o tiredness
C0015672|033|sensation of weakness
C0015672|033|decreased activity
C0015672|033|cannot finish adls
C0015672|033|decreased job performance
C0015672|033|not feeling rested
C0015672|033|persistent tiredness
C0015672|033|ongoing fatigue
C0015672|033|constant fatigue
C0015672|033|intermittent fatigue
C0015672|033|periodic fatigue
C0015672|033|worsening fatigue
C0015672|033|recurrent fatigue
C0015672|033|energy deficit
C0015672|033|vitality loss
C0015672|033|weakness
C0015672|033|generalized weakness
C0015672|033|focal weakness
C0015672|033|muscle weakness
C0015672|033|proximal weakness
C0015672|033|distal weakness
C0015672|033|asthenia
C0015672|033|paresis
C0015672|033|hemiparesis
C0015672|033|paraparesis
C0015672|033|quadriparesis
C0015672|033|tetraparesis
C0015672|033|myopathy
C0015672|033|fatigue
C0015672|033|malaise
C0015672|033|decreased strength
C0015672|033|low strength
C0015672|033|diminished strength
C0015672|033|loss of strength
C0015672|033|power loss
C0015672|033|reduced power
C0015672|033|motor deficit
C0015672|033|motor impairment
C0015672|033|flaccidity
C0015672|033|flaccid muscles
C0015672|033|muscular fatigue
C0015672|033|exertional fatigue
C0015672|033|neuromuscular weakness
C0015672|033|hyposthenia
C0015672|033|nm weakness
C0015672|033|decreased grip strength
C0015672|033|sluggish muscle response
C0015672|033|muscle atony
C0015672|033|muscle hypotonia
C0015672|033|floppy muscles
C0015672|033|muscle insufficiency
C0015672|033|myasthenia
C0015672|033|ppcm-related weakness
C0015672|033|cva-related weakness
C0015672|033|stroke-related weakness
C0015672|033|ischemic weakness
C0015672|033|nonischemic weakness
C0015672|033|chemo-induced weakness
C0015672|033|drug-induced weakness
C0015672|033|myocarditis-related weakness
C0015672|033|valvular-related weakness
C0015672|033|hypertensive weakness
C0015672|033|amyloid weakness
C0015672|033|tachycardia-induced weakness
C0015672|033|als-related weakness
C0015672|033|ms-related weakness
C0015672|033|parkinsonian weakness
C0015672|033|alcoholic weakness
C0015672|033|critical illness weakness
C0015672|033|periodic paralysis
C0015672|033|central weakness
C0015672|033|peripheral weakness
C0015672|033|monoparesis
C0015672|033|paresis rle
C0015672|033|paresis lle
C0015672|033|paresis rue
C0015672|033|paresis lue
C0015672|033|le weakness
C0015672|033|rle weakness
C0015672|033|lle weakness
C0015672|033|ue weakness
C0015672|033|rue weakness
C0015672|033|lue weakness
C0015672|033|diffuse weakness
C0015672|033|bilateral weakness
C0015672|033|unilateral weakness
C0015672|033|r-sided weakness
C0015672|033|l-sided weakness
C0015672|033|impaired muscle strength
C0015672|033|mobility impairment
C0015672|033|ambulatory weakness
C0015672|033|transient weakness
C0015672|033|chronic weakness
C0015672|033|acute weakness
C0015672|033|subjective weakness
C0015672|033|objective weakness
C0015672|033|myotonia
C0015672|033|em weakness
C0015672|033|functional weakness
C0015672|033|secondary weakness
C0015672|033|progressive weakness
C0015672|033|persistent weakness
C0015672|033|episodic weakness
C0015672|033|muscle deficit
C0015672|033|neuropathic weakness
C0015672|033|myopathic weakness
C0015672|033|limb weakness
C0015672|033|down-going strength
C0015672|033|paresis limb
C0015672|033|paresis extremity
C0015672|033|motor weakness
C0015672|033|loss of muscle function
C0015672|033|muscle deterioration
C0015672|033|muscle debility
C0015672|033|muscle flaccidity
C0015672|033|gait weakness
C0015672|033|muscle sluggishness
C0015672|033|frank weakness
C0015672|033|mild weakness
C0015672|033|moderate weakness
C0015672|033|marked weakness
C0015672|033|severe weakness
C0015672|033|pml-related weakness
C0015672|033|gbs-related weakness
C0015672|033|mnd weakness
C0015672|033|cidp-related weakness
C0015672|033|inflammatory weakness
C0015672|033|immune-mediated weakness
C0015672|033|cachectic weakness
C0015672|033|paraneoplastic weakness
C0015672|033|disuse weakness
C0015672|033|immobility-related weakness
C0015672|033|respiratory muscle weakness
C0015672|033|oculomotor weakness
C0015672|033|bulbar weakness
C0015672|033|facial weakness
C0015672|033|cranial nerve weakness
C0015672|033|truncal weakness
C0015672|033|core weakness
C0015672|033|hand weakness
C0015672|033|wrist drop
C0015672|033|foot drop
C0015672|033|muscle fatigability
C0015672|033|easy fatigability
C0015672|033|pem (post-exertional malaise)
C0015672|033|floppy baby
C0015672|033|motor neuron weakness
C0015672|033|neurogenic weakness
C0015672|033|recurrent weakness
C0015672|033|fluctuant weakness
C0015672|033|waxing/waning weakness
C0015672|033|emg-documented weakness
C0015672|033|exercise-induced weakness
C0015672|033|overuse weakness
C0015672|033|debilitation
C0015672|033|muscular debility
C0015672|033|myasthenic symptoms
C0015672|033|hypotonicity
C0015672|033|decreased tone
C0015672|033|drop attacks
C0015672|033|loss muscle bulk
C0015672|033|atrophic weakness
C0015672|033|lateralizing weakness
C0015672|033|symmetric weakness
C0015672|033|asymmetric weakness
C0015672|033|spastic weakness
C0015672|033|nonspastic weakness
C0015672|033|limb drift
C0015672|033|pronator drift
C0015672|033|clumsiness
C0015672|033|unsteady
C0015672|033|loss of antigravity strength
C0015672|033|muscle impairment
C0015672|033|poor muscle performance
C0015672|033|impaired performance
C0015672|033|decline muscle strength
C0015672|033|mechanical weakness
C0015672|033|myotoxicity
C0015672|033|toxic myopathy
C0015672|033|steroid-induced weakness
C0015672|033|corticosteroid myopathy
C0015672|033|paraplegic weakness
C0015672|033|plegic weakness
C0015672|033|flaccid paresis
C0015672|033|hypotonic weakness
C0015672|033|lower limb weakness
C0015672|033|upper limb weakness
C0015672|033|speech weakness
C0015672|033|dysarthric weakness
C0015672|033|pharyngeal weakness
C0015672|033|lingual weakness
C0015672|033|tongue weakness
C0015672|033|neck flexion weakness
C0015672|033|neck extension weakness
C0015672|033|axial weakness
C0015672|033|presynaptic weakness
C0015672|033|postsynaptic weakness
C0015672|033|distal limb weakness
C0015672|033|proximal limb weakness
C0015672|033|hand grip weakness
C0015672|033|paresis ues
C0015672|033|paresis les
C0015672|033|progressive myopathy
C0015672|033|myopathy nos
C0015672|033|myositis-related weakness
C0015672|033|limb heaviness
C0015672|033|heavy limbs
C0015672|033|muscle heaviness
C0015672|033|floppy infant
C0015672|033|myasthenic weakness
C0015672|033|neoplasm-related weakness
C0015672|033|critical illness myopathy
C0015672|033|systemic weakness
C0015672|033|pandysautonomia weakness
C5543391|033|low appetite
C5543391|033|↓ appetite
C5543391|033|decreased appetite
C5543391|033|dec appetite
C5543391|033|↓ po intake
C5543391|033|po intake ↓
C5543391|033|poor appetite
C5543391|033|reduced appetite
C5543391|033|loss of appetite
C5543391|033|appetite loss
C5543391|033|appetite ↓
C5543391|033|no appetite
C5543391|033|anorexia
C5543391|033|anorexic
C5543391|033|anorexia nervosa
C5543391|033|poor oral intake
C5543391|033|↓ oral intake
C5543391|033|low oral intake
C5543391|033|oral intake ↓
C5543391|033|diminished appetite
C5543391|033|diminished po intake
C5543391|033|appetite off
C5543391|033|avoiding food
C5543391|033|not eating well
C5543391|033|not eating
C5543391|033|decreased eating
C5543391|033|eating less
C5543391|033|appetite suppression
C5543391|033|anorexia (chemo-induced)
C5543391|033|chemo-induced anorexia
C5543391|033|chemo-induced appetite loss
C5543391|033|loss of appetite (chemo)
C5543391|033|appetite change
C5543391|033|poor po
C5543391|033|po poor
C5543391|033|s/p chemo ↓ appetite
C5543391|033|appetite poor
C5543391|033|low caloric intake
C5543391|033|↓ caloric intake
C5543391|033|hyporexia
C5543391|033|hyporexic
C5543391|033|poor feeding
C5543391|033|reduced feeding
C5543391|033|failure to thrive (ftt)
C5543391|033|ftt
C5543391|033|cachexia
C5543391|033|cancer cachexia
C5543391|033|tumor-induced anorexia
C5543391|033|nonischemic anorexia
C5543391|033|ischemic anorexia
C5543391|033|anorexia (myocarditis)
C5543391|033|tachycardia-induced anorexia
C5543391|033|myocarditis-related poor appetite
C5543391|033|chf-related loss of appetite
C5543391|033|valvular disease ↓ appetite
C5543391|033|appetite down
C5543391|033|poor intake
C5543391|033|decreased intake
C5543391|033|npo except meds
C5543391|033|intake less than baseline
C5543391|033|low nutritional intake
C5543391|033|food aversion
C5543391|033|feeding aversion
C5543391|033|reduced nutritional intake
C5543391|033|↓ interest in food
C5543391|033|reluctant to eat
C5543391|033|not hungry
C5543391|033|inappetent
C5543391|033|appetite suppressed
C5543391|033|self-restricted dietary intake
C5543391|033|poor nutrition
C5543391|033|voluntary starvation
C5543391|033|intentional anorexia
C5543391|033|starvation (anorexia)
C5543391|033|poor intake (ppcm)
C5543391|033|amyloidosis-related appetite loss
C5543391|033|amyloidosis poor appetite
C5543391|033|inadequate po intake
C5543391|033|low po
C5543391|033|low food consumption
C5543391|033|eating < normal
C5543391|033|intake < normal
C5543391|033|↓ food consumption
C5543391|033|diminished desire to eat
C5543391|033|unable to tolerate po
C5543391|033|appetite lacking
C5543391|033|decreased desire for food
C5543391|033|loss of interest in eating
C5543391|033|skipping meals
C5543391|033|refusing meals
C5543391|033|using appetite suppressants
C5543391|033|gi-related ↓ appetite
C5543391|033|hepatic anorexia
C5543391|033|heart failure anorexia
C5543391|033|cardiac cachexia
C5543391|033|ckd-related anorexia
C5543391|033|esrd-related poor appetite
C5543391|033|dialysis-related ↓ appetite
C5543391|033|uremic anorexia
C5543391|033|copd-related ↓ appetite
C5543391|033|hiv-related anorexia
C5543391|033|infection-related loss of appetite
C5543391|033|sepsis anorexia
C5543391|033|tb-related poor appetite
C5543391|033|anorexia secondary to disease
C5543391|033|malignancy-related ↓ appetite
C5543391|033|oncologic anorexia
C5543391|033|appetite complaint
C5543391|033|reduced caloric intake
C5543391|033|nutrition intake suboptimal
C5543391|033|nutrition: poor
C5543391|033|nutrition: decreased
C5543391|033|eats very little
C5543391|033|minimal po intake
C5543391|033|↓ consumption
C5543391|033|low dietary intake
C5543391|033|dietary intake reduced
C5543391|033|unable to eat
C5543391|033|feeding difficulty
C5543391|033|reluctance to feed
C5543391|033|anorexia (psychiatric)
C5543391|033|geriatric anorexia
C5543391|033|pediatric poor feeding
C5543391|033|hunger absent
C5543391|033|non-volitional ↓ intake
C5543391|033|self-limited po
C5543391|033|voluntarily not eating
C5543391|033|hypophagia
C5543391|033|hypophagic
C5543391|033|prn appetite loss
C5543391|033|drug-induced anorexia
C5543391|033|opioid-induced ↓ appetite
C5543391|033|antibiotic-induced ↓ appetite
C5543391|033|ssris - appetite loss
C5543391|033|steroid-induced ↓ appetite
C5543391|033|appetite suppressed (rx)
C5543391|033|stress-induced anorexia
C5543391|033|depression-related decreased appetite
C5543391|033|anxiety-related anorexia
C5543391|033|po intolerance
C5543391|033|unable to tolerate oral intake
C5543391|033|failure to eat
C5543391|033|refusal to eat
C5543391|033|appetite reduced
C5543391|033|appetite significantly ↓
C5543391|033|sarcopenia-related poor intake
C5543391|033|impaired appetite
C5543391|033|low feeding drive
C5543391|033|early satiety
C5543391|033|no desire for food
C5543391|033|satiety at low volumes
C5543391|033|perceived anorexia
C5543391|033|progressive decrease in appetite
C5543391|033|acute onset anorexia
C5543391|033|chronic poor appetite
C5543391|033|recurrent anorexia
C5543391|033|appetite disturbance
C5543391|033|low interest in food
C5543391|033|gastrointestinal symptoms - poor appetite
C5543391|033|post-op ↓ appetite
C5543391|033|post-infectious anorexia
C5543391|033|postpartum poor appetite
C5543391|033|pregnancy-related appetite loss
C5543391|033|appetite off since illness
C5543391|033|withdrew from eating
C5543391|033|low po tolerance
C5543391|033|poor caloric intake
C5543391|033|appetite not present
C5543391|033|cannot tolerate diet
C5543391|033|appetite declining
C5543391|033|eating reluctance
C5543391|033|no feeding
C5543391|033|neglecting meals
C5543391|033|adhf-related ↓ appetite
C5543391|033|low po desire
C5543391|033|lack of hunger
C5543391|033|reduced food preference
C5543391|033|reduced desire for food
C0003123|033|anorexia
C0003123|033|anorexic
C0003123|033|↓ appetite
C0003123|033|decreased appetite
C0003123|033|loss of appetite
C0003123|033|poor appetite
C0003123|033|reduced appetite
C0003123|033|anorexia nervosa
C0003123|033|cancer anorexia
C0003123|033|chemo-induced anorexia
C0003123|033|drug-induced anorexia
C0003123|033|appetite loss
C0003123|033|appetite suppression
C0003123|033|no appetite
C0003123|033|failure to eat
C0003123|033|refusing food
C0003123|033|not eating
C0003123|033|appetite reduction
C0003123|033|inappetence
C0003123|033|hyporexia
C0003123|033|appetite decline
C0003123|033|diminished appetite
C0003123|033|lack of appetite
C0003123|033|poor po intake
C0003123|033|anorexia-cachexia
C0003123|033|chf-related anorexia
C0003123|033|ckd-related anorexia
C0003123|033|esrd anorexia
C0003123|033|uremic anorexia
C0003123|033|gi-induced anorexia
C0003123|033|infectious anorexia
C0003123|033|psychogenic anorexia
C0003123|033|depression-related anorexia
C0003123|033|hepatic anorexia
C0003123|033|liver disease anorexia
C0003123|033|dementia anorexia
C0003123|033|dementia-related decreased appetite
C0003123|033|appetite off
C0003123|033|not interested in food
C0003123|033|patient not eating
C0003123|033|voluntary food restriction
C0003123|033|starvation
C0003123|033|no po
C0003123|033|↓ oral intake
C0003123|033|not tolerating po
C0003123|033|↓ food intake
C0003123|033|minimal intake
C0003123|033|reduced po intake
C0003123|033|decreased po
C0003123|033|refusal to eat
C0575081|033|gait abnormality
C0575081|033|abnormal gait
C0575081|033|gait disturbance
C0575081|033|abnormal gait pattern
C0575081|033|disordered gait
C0575081|033|ataxic gait
C0575081|033|gait ataxia
C0575081|033|unsteady gait
C0575081|033|walking difficulty
C0575081|033|disturbed ambulation
C0575081|033|abnormal ambulation
C0575081|033|ambulatory dysfunction
C0575081|033|abnormal walking
C0575081|033|impaired gait
C0575081|033|gait impairment
C0575081|033|ambulatory impairment
C0575081|033|difficulty walking
C0575081|033|impaired ambulation
C0575081|033|abnormal locomotion
C0575081|033|locomotor abnormality
C0575081|033|gait instability
C0575081|033|instability walking
C0575081|033|unstable gait
C0575081|033|gait dyspraxia
C0575081|033|shuffling gait
C0575081|033|festinating gait
C0575081|033|parkinsonian gait
C0575081|033|spastic gait
C0575081|033|spastic-ataxic gait
C0575081|033|hemiplegic gait
C0575081|033|hemiparetic gait
C0575081|033|diplegic gait
C0575081|033|scissoring gait
C0575081|033|scissor gait
C0575081|033|trendelenburg gait
C0575081|033|waddling gait
C0575081|033|cerebellar gait
C0575081|033|sensory ataxia
C0575081|033|apraxic gait
C0575081|033|myopathic gait
C0575081|033|steppage gait
C0575081|033|neuropathic gait
C0575081|033|foot drop gait
C0575081|033|paraparetic gait
C0575081|033|high-stepping gait
C0575081|033|magnetic gait
C0575081|033|hypokinetic gait
C0575081|033|bradykinetic gait
C0575081|033|tabetic gait
C0575081|033|choreiform gait
C0575081|033|antalgic gait
C0575081|033|limping gait
C0575081|033|walking abnormality
C0575081|033|walking disturbance
C0575081|033|abnl gait
C0575081|033|gait abnl
C0575081|033|gait dis
C0575081|033|gait dist
C0575081|033|impaired walking
C0575081|033|mobility impairment
C0575081|033|mobility abnormality
C0575081|033|decreased mobility
C0575081|033|gait dysfunction
C0575081|033|gait unsteadiness
C0575081|033|wide-based gait
C0575081|033|narrow-based gait
C0575081|033|small steps gait
C0575081|033|short stride gait
C0575081|033|gait freezing
C0575081|033|gait block
C0575081|033|propulsive gait
C0575081|033|paretic gait
C0575081|033|staggering gait
C0575081|033|drunken gait
C0575081|033|elderly gait disturbance
C0575081|033|frontal gait disorder
C0575081|033|gait disorder nos
C0575081|033|abnormal gait nos
C0575081|033|gait disturbance nos
C0575081|033|difficulty ambulating
C0575081|033|impaired gross mobility
C0575081|033|slow gait
C0575081|033|slowness walking
C0575081|033|gait slowness
C0575081|033|cautious gait
C0575081|033|gait hesitation
C0575081|033|equinus gait
C0575081|033|toe-walking
C0575081|033|toe gait
C0575081|033|calcaneal gait
C0575081|033|heel-walking
C0575081|033|clumsy gait
C0575081|033|abnl ambulation
C0575081|033|ms-related gait dysfunction
C0575081|033|parkinson's gait
C0575081|033|hemiplegic walking
C0575081|033|functional gait disorder
C0575081|033|conversion gait
C0575081|033|psychogenic gait
C0575081|033|malingered gait
C0575081|033|tremor during gait
C0575081|033|dystonic gait
C0575081|033|spastic-hemiplegic gait
C0575081|033|flaccid gait
C0575081|033|choreaform gait
C0575081|033|basal ganglia gait disorder
C0575081|033|extrapyramidal gait disorder
C0575081|033|gait apraxia
C0575081|033|gait difficulty
C0575081|033|abnormal stride
C0575081|033|gait deviation
C0575081|033|gait change
C0575081|033|gait deficit
C0575081|033|poor gait
C0575081|033|altered gait
C0575081|033|altered ambulation
C0575081|033|disrupted gait
C0575081|033|gait impairment due to stroke
C0575081|033|post-stroke gait
C0575081|033|ischemic gait abnormality
C0575081|033|chemo-induced gait abnormality
C0575081|033|myelopathy-related gait disorder
C0575081|033|radiculopathy gait abnormality
C0575081|033|als-related gait abnormality
C0575081|033|motor neuron gait deficit
C0575081|033|pyramidal gait
C0575081|033|spinal gait disturbance
C0575081|033|cerebral palsy gait
C0575081|033|cp gait
C0575081|033|demyelinating gait
C0575081|033|peripheral neuropathy gait
C0575081|033|diabetic gait disturbance
C0575081|033|amyloid gait abnormality
C0575081|033|hypertensive gait disorder
C0575081|033|valvular gait disorder
C0575081|033|tachycardia-induced gait abnormality
C0575081|033|ppcm gait abnormality
C0575081|033|myocarditis gait abnormality
C0575081|033|mixed pattern gait
C0575081|033|sensory-motor gait disturbance
C0575081|033|posterior column gait disorder
C0575081|033|spastic-paraparetic gait
C0575081|033|bilateral gait disturbance
C0575081|033|bilateral leg gait abnormality
C0575081|033|spastic quadriparetic gait
C0575081|033|quadriparetic gait
C0575081|033|unmotivated gait
C0575081|033|weak gait
C0575081|033|loss of gait automation
C0575081|033|frontal ataxia
C0575081|033|subcortical gait disturbance
C0575081|033|akinetic gait
C0575081|033|hypometric gait
C0575081|033|dyskinetic gait
C0575081|033|hyperkinetic gait
C0575081|033|swaying gait
C0575081|033|leaning gait
C0575081|033|lateralized gait
C0575081|033|ill-compensated gait
C0575081|033|postural gait abnormality
C0575081|033|drop foot gait
C0575081|033|hemiparetic walking
C0575081|033|toe drag gait
C0575081|033|step-page gait
C0575081|033|stooped gait
C0575081|033|stiff-legged gait
C0575081|033|genu recurvatum gait
C0575081|033|myotonic gait
C0575081|033|ataxia
C0575081|033|gmf dysfunction
C0575081|033|gmf deficit
C0575081|033|trendelenburg sign
C0575081|033|incoordinated gait
C0575081|033|nonphysiologic gait
C0575081|033|friction gait
C0575081|033|gait deviation due to spasticity
C0575081|033|spasticity-related gait change
C0575081|033|spastic diplegic gait
C0575081|033|dysfunctional stride
C0575081|033|gait variance
C0241981|033|impaired balance
C0241981|033|balance impairment
C0241981|033|unsteady gait
C0241981|033|gait instability
C0241981|033|ataxia
C0241981|033|vestibular dysfunction
C0241981|033|loss of balance
C0241981|033|postural instability
C0241981|033|impaired coordination
C0241981|033|equilibrium disturbance
C0241981|033|gait disturbance
C0241981|033|unsteadiness
C0241981|033|dizziness
C0241981|033|disequilibrium
C0241981|033|vertigo
C0241981|033|unsteady on feet
C0241981|033|wobbling gait
C0241981|033|staggering
C0241981|033|romberg positive
C0241981|033|wide-based gait
C0241981|033|abnormal gait
C0241981|033|waddling gait
C0241981|033|lurching gait
C0241981|033|drunken gait
C0241981|033|gait ataxia
C0241981|033|impaired proprioception
C0241981|033|impaired vestibular function
C0241981|033|labyrinthine dysfunction
C0241981|033|cerebellar ataxia
C0241981|033|sensory ataxia
C0241981|033|vestibular ataxia
C0241981|033|spinocerebellar ataxia
C0241981|033|paraparesis
C0241981|033|spastic gait
C0241981|033|toe-walking
C0241981|033|impairment of equilibrium
C0241981|033|impaired stance
C0241981|033|swaying
C0241981|033|gait abnormality
C0241981|033|shuffling gait
C0241981|033|parkinsonian gait
C0241981|033|gait deviation
C0241981|033|sway-positive
C0241981|033|antalgic gait
C0241981|033|hemiparetic gait
C0241981|033|ataxic gait
C0241981|033|impaired ambulation
C0241981|033|poor balance
C0241981|033|abnormal tandem gait
C0241981|033|abnormal heel-to-toe walk
C0241981|033|impaired tandem gait
C0241981|033|instability
C0241981|033|gait disorder
C0241981|033|gait unsteadiness
C0241981|033|marching unsteadily
C0241981|033|perceived imbalance
C0241981|033|oscillopsia
C0241981|033|feelings of imbalance
C0241981|033|impaired postural control
C0241981|033|abnormal posture
C0241981|033|bilateral leg unsteadiness
C0241981|033|loss of proprioception
C0241981|033|falling tendencies
C0241981|033|near falls
C0241981|033|off-balance
C0241981|033|loss of stability
C0241981|033|gait uncoordination
C0241981|033|drifting to side
C0241981|033|proprioceptive deficit
C0241981|033|sway on standing
C0241981|033|impaired romberg
C0241981|033|positive romberg
C0241981|033|disordered equilibrium
C0241981|033|gait dyspraxia
C0241981|033|dysmetria
C0241981|033|dysequilibrium
C0241981|033|locomotor ataxia
C0241981|033|veering
C0241981|033|poor righting reflex
C0241981|033|abnormal righting response
C0241981|033|truncal ataxia
C0241981|033|hypotonic gait
C0241981|033|gait freezing
C0241981|033|festination
C0241981|033|drop attacks
C0241981|033|frequent stumbles
C0241981|033|frequent falls
C0241981|033|abnormal gait mechanics
C0241981|033|limb incoordination
C0241981|033|balance deficit
C0241981|033|balance disorder
C0241981|033|compromised balance
C0241981|033|equilibrium disorder
C0241981|033|abnormal balance
C0241981|033|impaired verticality
C0241981|033|standing instability
C0241981|033|abnormal balance test
C0241981|033|proprioceptive gait disorder
C0241981|033|myopathy gait
C0241981|033|neuropathic gait
C0241981|033|steppage gait
C0241981|033|acute vestibulopathy
C0241981|033|central vestibulopathy
C0241981|033|peripheral vestibulopathy
C0241981|033|cerebellopathy
C0241981|033|ischemic ataxia
C0241981|033|nonischemic ataxia
C0241981|033|stroke-related instability
C0241981|033|tbi-related balance loss
C0241981|033|cva with gait disturbance
C0241981|033|ms-related ataxia
C0241981|033|parkinson’s gait disturbance
C0241981|033|chemo-induced ataxia
C0241981|033|medication-induced imbalance
C0241981|033|alcohol-induced ataxia
C0241981|033|diabetic ataxia
C0241981|033|amyloid neuropathy gait
C0241981|033|thiamine-deficient ataxia
C0241981|033|vitamin b12 deficiency gait
C0241981|033|myelopathy-induced gait impairment
C0241981|033|spinal stenosis–related balance loss
C0241981|033|peripheral neuropathy–related imbalance
C0241981|033|sensory neuropathy gait
C0241981|033|tachycardia-induced syncope with falls
C0241981|033|ppcm-related unsteady gait
C0241981|033|chf with instability
C0241981|033|hypertensive encephalopathy ataxia
C0241981|033|cerebellar infarct with imbalance
C0241981|033|vertebrobasilar insufficiency with ataxia
C0241981|033|valvular disease with falls
C0241981|033|meniere’s disease imbalance
C0241981|033|bppv imbalance
C0241981|033|ototoxicity with gait disturbance
C0241981|033|presbystasis
C0241981|033|areflexia with unsteady gait
C0241981|033|ortho hypotension with falls
C0241981|033|acute labyrinthitis
C0241981|033|chronic imbalance
C0241981|033|idiopathic ataxia
C0241981|033|post-ictal unsteadiness
C0241981|033|post-surgical imbalance
C0241981|033|age-related imbalance
C0241981|033|impaired walk
C0241981|033|coordination deficit
C0241981|033|uncoordinated gait
C0241981|033|disordered gait
C0241981|033|impaired locomotion
C0241981|033|impaired walking stability
C0241981|033|tripping easily
C0241981|033|impaired stance control
C0241981|033|marked gait disturbance
C0241981|033|walks with assistance
C0241981|033|requires mobility aid
C0241981|033|frequent wall walking
C0241981|033|unstable gait
C0241981|033|instability on ambulation
C0241981|033|poor postural stability
C0241981|033|unsteady when turning
C0241981|033|unsteady standing
C0241981|033|poor dynamic balance
C0241981|033|deficient balance response
C0241981|033|impaired dynamic equilibrium
C0241981|033|imbalance
C0241981|033|bos-wide gait
C0241981|033|need for assistive device due to balance
C0241981|033|use of cane for balance
C1405979|033|radiation necrosis
C1405979|033|radiation-induced necrosis
C1405979|033|post-radiation necrosis
C1405979|033|postirradiation necrosis
C1405979|033|radionecrosis
C1405979|033|radiation-related necrosis
C1405979|033|rt necrosis
C1405979|033|radio-necrosis
C1405979|033|irradiation necrosis
C1405979|033|necrosis secondary to radiation
C1405979|033|necrosis d/t radiation
C1405979|033|necrosis s/p radiation
C1405979|033|necrosis d/t rt
C1405979|033|necrosis s/p rt
C1405979|033|necrosis s/p irradiation
C1405979|033|post-radiotherapy necrosis
C1405979|033|radiotherapy necrosis
C1405979|033|necrosis following ionizing radiation
C1405979|033|ionizing radiation necrosis
C1405979|033|necrosis due to radiotherapy
C1405979|033|post-rt necrosis
C1405979|033|radiation necrotic changes
C1405979|033|radionecrotic lesion
C1405979|033|radiation injury with necrosis
C1405979|033|radiation effect necrosis
C1405979|033|secondary radiation necrosis
C1405979|033|delayed radiation necrosis
C1405979|033|delayed radionecrosis
C1405979|033|late rt necrosis
C1405979|033|late radiation necrosis
C1405979|033|chronic radiation necrosis
C1405979|033|chronic radionecrosis
C1405979|033|focal radiation necrosis
C1405979|033|multifocal radiation necrosis
C1405979|033|gliocentric radiation necrosis
C1405979|033|nonischemic radiation necrosis
C1405979|033|ischemic radiation necrosis
C1405979|033|necrosis due to therapeutic irradiation
C1405979|033|therapy-induced necrosis
C1405979|033|treatment-induced necrosis
C1405979|033|necrosis post-external beam rt
C1405979|033|necrosis secondary to ebrt
C1405979|033|ebrt necrosis
C1405979|033|gamma knife necrosis
C1405979|033|stereotactic radiosurgery necrosis
C1405979|033|srs necrosis
C1405979|033|srt necrosis
C1405979|033|sbrt necrosis
C1405979|033|cns radiation necrosis
C1405979|033|brain radiation necrosis
C1405979|033|cerebral radiation necrosis
C1405979|033|myocardial radiation necrosis
C1405979|033|hepatic radiation necrosis
C1405979|033|pancreatic radiation necrosis
C1405979|033|soft tissue radiation necrosis
C1405979|033|cutaneous radiation necrosis
C1405979|033|skin radiation necrosis
C1405979|033|lung radiation necrosis
C1405979|033|pulmonary radiation necrosis
C1405979|033|bone radiation necrosis
C1405979|033|mandibular radiation necrosis
C1405979|033|mandibular radionecrosis
C1405979|033|osteoradionecrosis
C1405979|033|radionecrosis of bone
C1405979|033|radionecrosis jaw
C1405979|033|radiation-induced bone necrosis
C1405979|033|soft tissue radionecrosis
C1405979|033|necrosis from rt
C1405979|033|necrosis from srs
C1405979|033|necrosis from radiosurgery
C1405979|033|necrosis from sbrt
C1405979|033|necrosis from gamma knife
C1405979|033|post-radiation necrotic change
C1405979|033|necrosis after irradiation
C1405979|033|necrosis following radiation therapy
C1405979|033|necrosis 2/2 radiation
C1405979|033|d/t rt necrosis
C1405979|033|post-xrt necrosis
C1405979|033|xrt necrosis
C1405979|033|ir necrosis
C1405979|033|necrosis s/p xrt
C1405979|033|necrosis d/t xrt
C1405979|033|necrosis post-xrt
C1405979|033|necrosis related to irradiation
C1405979|033|necrosis associated with radiation
C1405979|033|radiation damage with necrosis
C1405979|033|radiation-induced tissue necrosis
C1405979|033|tissue radionecrosis
C1405979|033|necrosis secondary to radiotherapy
C1405979|033|post-irradiation necrosis
C1405979|033|necrosis after beam therapy
C1405979|033|tissue death due to rt
C1405979|033|necrosis from therapeutic irradiation
C1405979|033|post-treatment necrosis (radiation)
C1405979|033|postradiosurgical necrosis
C1405979|033|sbrt-related necrosis
C1405979|033|srt-related necrosis
C1405979|033|stereotactic rt necrosis
C1405979|033|post-gamma knife necrosis
C1405979|033|gamma knife-induced necrosis
C1405979|033|irradiation effect necrosis
C1405979|033|irradiation-related necrosis
C1405979|033|necrosis subsequent to radiation
C1405979|033|necrosis subsequent to rt
C1405979|033|necrosis post radiotherapy
C1405979|033|necrosis after rt
C1405979|033|irradiation-associated necrosis
C1392786|033|cognitive dysfunction
C1392786|033|cognitive impairment
C1392786|033|cognitive decline
C1392786|033|cognitive deficits
C1392786|033|cognitive disturbance
C1392786|033|cognition impaired
C1392786|033|cognition changes
C1392786|033|altered cognition
C1392786|033|memory loss
C1392786|033|memory impairment
C1392786|033|forgetfulness
C1392786|033|short-term memory loss
C1392786|033|long-term memory loss
C1392786|033|confusion
C1392786|033|disorientation
C1392786|033|altered mental status
C1392786|033|ams
C1392786|033|encephalopathy
C1392786|033|delirium
C1392786|033|delirious
C1392786|033|acute mental status change
C1392786|033|fluctuating mental status
C1392786|033|clouded mentation
C1392786|033|mentation changes
C1392786|033|slowed mentation
C1392786|033|impaired executive function
C1392786|033|executive dysfunction
C1392786|033|difficulty concentrating
C1392786|033|concentration deficit
C1392786|033|decreased attention span
C1392786|033|attention deficit
C1392786|033|inattention
C1392786|033|impaired attention
C1392786|033|poor recall
C1392786|033|impaired recall
C1392786|033|impaired judgment
C1392786|033|judgment deficits
C1392786|033|difficulty making decisions
C1392786|033|reversible cognitive impairment
C1392786|033|irreversible cognitive impairment
C1392786|033|mild cognitive impairment
C1392786|033|mci
C1392786|033|dementia
C1392786|033|demented
C1392786|033|early-onset dementia
C1392786|033|late-onset dementia
C1392786|033|progressive cognitive decline
C1392786|033|vascular cognitive impairment
C1392786|033|ischemic cognitive impairment
C1392786|033|ischemic encephalopathy
C1392786|033|post-stroke cognitive changes
C1392786|033|stroke-related cognitive decline
C1392786|033|non-ischemic cognitive changes
C1392786|033|hypoxic encephalopathy
C1392786|033|hypoxic cognitive dysfunction
C1392786|033|chemo brain
C1392786|033|chemo-induced cognitive changes
C1392786|033|chemo-related cognitive impairment
C1392786|033|tumor-related cognitive change
C1392786|033|brain metastases cognitive effect
C1392786|033|radiation-induced cognitive decline
C1392786|033|amyloid-related cognitive impairment
C1392786|033|alzheimer's type changes
C1392786|033|ad-type dementia
C1392786|033|frontotemporal cognitive impairment
C1392786|033|lewy body cognitive dysfunction
C1392786|033|parkinson's-related cognitive change
C1392786|033|pd dementia
C1392786|033|ath-related cognitive dysfunction
C1392786|033|atherosclerotic cognitive impairment
C1392786|033|hypertensive encephalopathy
C1392786|033|hypertensive cognitive decline
C1392786|033|metabolic encephalopathy
C1392786|033|hepatic encephalopathy
C1392786|033|uremic encephalopathy
C1392786|033|sepsis-associated encephalopathy
C1392786|033|toxic-metabolic encephalopathy
C1392786|033|medication-related cognitive impairment
C1392786|033|polypharmacy-induced cognitive change
C1392786|033|sedative-induced confusion
C1392786|033|delirium due to meds
C1392786|033|alcohol-related cognitive dysfunction
C1392786|033|wernicke's encephalopathy
C1392786|033|korsakoff psychosis
C1392786|033|post-ictal confusion
C1392786|033|postictal cognitive changes
C1392786|033|epileptic cognitive dysfunction
C1392786|033|autoimmune encephalopathy
C1392786|033|paraneoplastic encephalopathy
C1392786|033|infectious encephalopathy
C1392786|033|hiv-associated neurocognitive disorder
C1392786|033|neurocognitive disorder
C1392786|033|mild neurocognitive disorder
C1392786|033|major neurocognitive disorder
C1392786|033|cns dysfunction
C1392786|033|brain fog
C1392786|033|slowed cognition
C1392786|033|mental slowing
C1392786|033|mental clouding
C1392786|033|diminished cognition
C1392786|033|reduced cognitive capacity
C1392786|033|task management difficulty
C1392786|033|slowed thought process
C1392786|033|impaired thought process
C1392786|033|slowed reaction time
C1392786|033|reduced mental clarity
C1392786|033|mental dullness
C1392786|033|cognitive slowing
C1392786|033|depressive pseudodementia
C1392786|033|mood-related cognitive dysfunction
C1392786|033|psychosis-related cognitive change
C1392786|033|schizophrenia cognitive deficits
C1392786|033|bipolar cognitive dysfunction
C1392786|033|anoxic encephalopathy
C1392786|033|co poisoning cognitive effect
C1392786|033|encephalopathic
C1392786|033|icu psychosis
C1392786|033|hospital-acquired delirium
C1392786|033|postoperative cognitive dysfunction
C1392786|033|sundowning
C1392786|033|pre-dementia state
C1392786|033|prodromal dementia
C1392786|033|subcortical dementia
C1392786|033|cortical dementia
C1392786|033|microvascular cognitive impairment
C1392786|033|subcortical ischemic cognitive change
C1392786|033|tbi cognitive deficits
C1392786|033|concussion cognitive changes
C1392786|033|blast injury cognitive change
C1392786|033|chronic traumatic encephalopathy
C1392786|033|huntington's cognitive impairment
C1392786|033|huntington's dementia
C1392786|033|wilson's disease cognitive change
C1392786|033|lyme neuroborreliosis cognitive effect
C1392786|033|post-covid cognitive dysfunction
C1392786|033|covid brain fog
C1392786|033|pasc cognitive change
C1392786|033|fatigue-related cognitive impairment
C1392786|033|sleep deprivation cognitive deficits
C1392786|033|obstructive sleep apnea cognitive change
C1392786|033|osa cognitive impairment
C1392786|033|drug-induced cognitive dysfunction
C1392786|033|thc-related cognitive change
C1392786|033|opioid-associated cognition change
C1392786|033|polytrauma cognitive deficits
C1392786|033|emotional distress-related cognition change
C1392786|033|adjustment disorder with cognitive symptoms
C1392786|033|adolescent cognitive changes
C1392786|033|geriatric cognitive decline
C1392786|033|aging-related cognitive change
C1392786|033|senile dementia
C1392786|033|senile cognitive changes
C1392786|033|mci-amnestic
C1392786|033|mci-nonamnestic
C1392786|033|attention/executive dysfunction
C1392786|033|language dysfunction
C1392786|033|praxis impairment
C1392786|033|visuospatial dysfunction
C1392786|033|agitation with cognitive impairment
C1392786|033|wandering with cognitive disorder
C1392786|033|anosognosia
C1392786|033|aphasia with cognitive decline
C1392786|033|agraphia/cognitive changes
C1392786|033|alexia/cognitive issues
C1392786|033|dysexecutive syndrome
C1392786|033|multifactorial cognitive impairment
C1392786|033|delirium superimposed on dementia
C0011206|033|delirium
C0011206|033|acute confusional state
C0011206|033|acs
C0011206|033|icu delirium
C0011206|033|hospital-acquired delirium
C0011206|033|acute brain failure
C0011206|033|subsyndromal delirium
C0011206|033|hyperactive delirium
C0011206|033|hypoactive delirium
C0011206|033|mixed delirium
C0011206|033|postoperative delirium
C0011206|033|post-op delirium
C0011206|033|post-anesthesia delirium
C0011206|033|emergence delirium
C0011206|033|agitated delirium
C0011206|033|toxic delirium
C0011206|033|metabolic delirium
C0011206|033|hepatic encephalopathy
C0011206|033|septic encephalopathy
C0011206|033|infectious delirium
C0011206|033|alcohol withdrawal delirium
C0011206|033|delirium tremens
C0011206|033|benzodiazepine withdrawal delirium
C0011206|033|drug-induced delirium
C0011206|033|chemo-induced delirium
C0011206|033|medication-induced delirium
C0011206|033|iatrogenic delirium
C0011206|033|icu psychosis
C0011206|033|sun-downing
C0011206|033|sundowning syndrome
C0011206|033|sundown syndrome
C0011206|033|acute encephalopathy
C0011206|033|fluctuating mental status
C0011206|033|waxing-waning mental status
C0011206|033|altered mental status
C0011206|033|ams
C0011206|033|mental status changes
C0011206|033|acute ams
C0011206|033|encephalopathic changes
C0011206|033|paranoid delirium
C0011206|033|delirious state
C0011206|033|clouded sensorium
C0011206|033|acute organic brain syndrome
C0011206|033|confusional syndrome
C0011206|033|toxic confusional state
C0011206|033|postictal confusion
C0011206|033|delirium superimposed on dementia
C0011206|033|delirium-on-dementia
C0011206|033|delirium of mixed etiology
C0011206|033|covid delirium
C0011206|033|hypoxemic delirium
C0011206|033|urosepsis delirium
C0011206|033|sepsis-associated delirium
C0011206|033|delirium due to uti
C0011206|033|delirium due to pneumonia
C0011206|033|perceptual disturbance
C0011206|033|psychomotor agitation
C0011206|033|psychomotor disturbance
C0011206|033|transient cognitive impairment
C0011206|033|transient delirium
C0011206|033|acute psychosis (delirium type)
C0011206|033|agitated confusion
C0011206|033|disorganized thinking
C0011206|033|attention deficit (acute)
C0011206|033|acute cognitive dysfunction
C0011206|033|perioperative delirium
C0011206|033|delirium of elderly
C0011206|033|delirium in dementia
C0011206|033|terminal delirium
C0011206|033|end-of-life delirium
C0011206|033|delirium in palliative care
C0011206|033|uremic encephalopathy
C0011206|033|hepatic delirium
C0011206|033|delirium secondary to infection
C0011206|033|delirium secondary to metabolic encephalopathy
C0011206|033|nonconvulsive status epilepticus with confusional state
C0011206|033|post-cardiac surgery delirium
C0011206|033|trauma-related delirium
C0011206|033|withdrawal delirium
C0011206|033|anticholinergic toxicity
C0011206|033|anticholinergic delirium
C0011206|033|delirium due to medication
C0011206|033|cns toxicity (delirium)
C0011206|033|delirium state
C0011206|033|delirium episode
C0011206|033|acute onset confusion
C0011206|033|delirious episode
C0011206|033|confusional episode
C0011206|033|acute cognitive change
C0011206|033|acute mental status change
C0011206|033|catatonic delirium
C0011206|033|poststroke delirium
C0011206|033|delirium due to stroke
C0011206|033|opiate-induced delirium
C0011206|033|pain control delirium
C0011206|033|cardiac surgery delirium
C0011206|033|anoxic delirium
C0011206|033|sleep deprivation delirium
C0011206|033|encephalopathic delirium
C0011206|033|toxic-metabolic encephalopathy
C0011206|033|endocrine delirium
C0011206|033|thyrotoxic encephalopathy
C0011206|033|thyroid storm delirium
C0011206|033|delirium due to cerebral hypoperfusion
C0011206|033|pediatric delirium
C0011206|033|delirium in children
C0011206|033|hepatic failure delirium
C0011206|033|delirium due to renal failure
C0011206|033|reversible encephalopathy
C0011206|033|wernicke's encephalopathy
C0011206|033|alcohol-related delirium
C0011206|033|stimulant-induced delirium
C0011206|033|delirium nos
C0011206|033|acute delirium episode
C0011206|033|delirium of advanced age
C0011206|033|delirium of critical illness
C0011206|033|delirium by dsm criteria
C0497327|033|dementia
C0497327|033|demented
C0497327|033|major neurocognitive disorder
C0497327|033|chronic cognitive impairment
C0497327|033|cognitive decline
C0497327|033|cognitive dysfunction
C0497327|033|memory loss syndrome
C0497327|033|progressive cognitive decline
C0497327|033|senile dementia
C0497327|033|senile dem
C0497327|033|senile degeneration
C0497327|033|senile brain disease
C0497327|033|presenile dementia
C0497327|033|vascular dementia
C0497327|033|multi-infarct dementia
C0497327|033|arteriosclerotic dementia
C0497327|033|ischemic dementia
C0497327|033|post-stroke dementia
C0497327|033|alzheimer disease
C0497327|033|ad
C0497327|033|alzheimer's dementia
C0497327|033|alzheimer-type dementia
C0497327|033|mixed dementia
C0497327|033|dementia with lewy bodies
C0497327|033|lewy body dementia
C0497327|033|frontotemporal dementia
C0497327|033|pick disease
C0497327|033|pick's dementia
C0497327|033|subcortical dementia
C0497327|033|huntington dementia
C0497327|033|huntington's dementia
C0497327|033|hd dementia
C0497327|033|parkinsonian dementia
C0497327|033|parkinson's dementia
C0497327|033|parkinsonism with dementia
C0497327|033|alcoholic dementia
C0497327|033|wernicke-korsakoff syndrome
C0497327|033|hiv-associated dementia
C0497327|033|aids-dementia complex
C0497327|033|hiv dementia
C0497327|033|posttraumatic dementia
C0497327|033|traumatic dementia
C0497327|033|tbi-related dementia
C0497327|033|chronic traumatic encephalopathy
C0497327|033|creutzfeldt-jakob dementia
C0497327|033|creutzfeldt-jakob disease
C0497327|033|prion dementia
C0497327|033|rapidly progressive dementia
C0497327|033|amyloid dementia
C0497327|033|autoimmune dementia
C0497327|033|hashimoto encephalopathy
C0497327|033|he dementia
C0497327|033|normal pressure hydrocephalus dementia
C0497327|033|nph dementia
C0497327|033|hydrocephalic dementia
C0497327|033|hepatic encephalopathy with dementia
C0497327|033|liver-related dementia
C0497327|033|hepatic dementia
C0497327|033|dialysis dementia
C0497327|033|uremic dementia
C0497327|033|metabolic dementia
C0497327|033|toxic dementia
C0497327|033|chemo-induced dementia
C0497327|033|chemotherapy-related cognitive impairment
C0497327|033|paraneoplastic dementia
C0497327|033|hypoxic-ischemic encephalopathy with dementia
C0497327|033|hie dementia
C0497327|033|hypoxic-ischemic dementia
C0497327|033|postanoxic dementia
C0497327|033|hypoglycemic dementia
C0497327|033|endocrine dementia
C0497327|033|thyroid dementia
C0497327|033|thyroid-related cognitive impairment
C0497327|033|syphilitic dementia
C0497327|033|neurosyphilis with dementia
C0497327|033|progressive paralytic dementia
C0497327|033|progressive general paralysis of the insane
C0497327|033|dementia praecox
C0497327|033|madness
C0497327|033|organic brain syndrome
C0497327|033|chronic organic brain disorder
C0497327|033|cerebral degeneration
C0497327|033|brain failure
C0497327|033|global cognitive dysfunction
C0497327|033|general cognitive decline
C0497327|033|chronic encephalopathy
C0497327|033|irreversible cognitive decline
C0497327|033|idiopathic dementia
C0497327|033|primary dementia
C0497327|033|secondary dementia
C0497327|033|drug-induced cognitive impairment
C0497327|033|iatrogenic dementia
C0497327|033|nos dementia
C0497327|033|not otherwise specified dementia
C0497327|033|late-onset dementia
C0497327|033|early-onset dementia
C0497327|033|juvenile dementia
C0497327|033|mild dementia
C0497327|033|moderate dementia
C0497327|033|severe dementia
C0497327|033|advanced dementia
C0497327|033|terminal dementia
C0497327|033|rapid-onset dementia
C0497327|033|progressive dementia
C0497327|033|static dementia
C0497327|033|potentially reversible dementia
C0497327|033|irreversible dementia
C0497327|033|prodromal dementia
C0497327|033|amnestic syndrome
C0497327|033|amnestic disorder
C0497327|033|korsakoff dementia
C0497327|033|wernicke dementia
C0497327|033|non-ad dementia
C0497327|033|non-alzheimer dementia
C0497327|033|prion-related dementia
C0497327|033|motor neuron disease dementia
C0497327|033|als dementia
C0497327|033|amyotrophic lateral sclerosis dementia
C0497327|033|peripheral neuropathy with dementia
C0497327|033|diffuse lewy body disease
C0497327|033|familial dementia
C0497327|033|inherited dementia
C0497327|033|cerebral amyloid angiopathy-related dementia
C0497327|033|caa dementia
C0497327|033|cadasil-related dementia
C0497327|033|cadasil dementia
C0497327|033|notch3 dementia
C0497327|033|binswanger disease
C0497327|033|binswanger's dementia
C0497327|033|subcortical arteriosclerotic encephalopathy
C0497327|033|reversible dementia
C0497327|033|parkinson-plus dementia
C0497327|033|progressive supranuclear palsy dementia
C0497327|033|psp dementia
C0497327|033|corticobasal degeneration dementia
C0497327|033|cbd dementia
C0497327|033|dementia syndrome
C0497327|033|aphasic dementia
C0497327|033|semantic dementia
C0497327|033|logopenic dementia
C0497327|033|primary progressive aphasia
C0497327|033|behavioral variant ftd
C0497327|033|semantic variant ppa
C0497327|033|nonfluent variant ppa
C0497327|033|nph cognitive impairment
C0497327|033|postinfectious dementia
C0497327|033|postmeningitic dementia
C0497327|033|herpes simplex encephalitis with dementia
C0497327|033|autoimmune encephalitis with dementia
C0497327|033|syndrome of dementia
C0497327|033|dementia-like syndrome
C0497327|033|mild cognitive impairment progressing to dementia
C0497327|033|mci progressing to dementia
C0497327|033|mci-to-dementia
C0497327|033|major ncd
C0497327|033|progressive memory loss
C0497327|033|intellectual deterioration
C0497327|033|generalized cognitive impairment
C0021125|033|impulsivity
C0021125|033|impulsive tendencies
C0021125|033|impulse control deficit
C0021125|033|impaired impulse control
C0021125|033|disinhibition
C0021125|033|disinhibited behavior
C0021125|033|behavioral disinhibition
C0021125|033|poor impulse control
C0021125|033|difficulty controlling impulses
C0021125|033|loss of impulse control
C0021125|033|acting on impulse
C0021125|033|compulsive urges
C0021125|033|compulsive actions
C0021125|033|lack of inhibition
C0021125|033|lack of self-control
C0021125|033|difficulty delaying gratification
C0021125|033|acts without thinking
C0021125|033|rash behavior
C0021125|033|impulsive acts
C0021125|033|impulsive responding
C0021125|033|impulsive actions
C0021125|033|impaired behavioral regulation
C0021125|033|reduced impulse control
C0021125|033|frontal lobe disinhibition
C0021125|033|frontal release
C0021125|033|auto-impulsive behavior
C0021125|033|impulsive decision-making
C0021125|033|poor behavioral inhibition
C0021125|033|diminished impulse control
C0021125|033|unrestrained behavior
C0021125|033|uncontrolled impulses
C0021125|033|lack of self-restraint
C0021125|033|executive dysfunction—impulsivity
C0021125|033|prefrontal syndrome—impulsivity
C0021125|033|hyperactivity—impulsivity
C0021125|033|bid (behavioral impulse dysregulation)
C0021125|033|icd (impulse control disorder)
C0021125|033|adhd-impulsivity
C0021125|033|addictive behavior
C0021125|033|mania—impulsivity
C0021125|033|manic impulsivity
C0021125|033|bpad—impulsivity
C0021125|033|tbi—disinhibition
C0021125|033|post-stroke impulsivity
C0021125|033|ischemic-frontal impulsivity
C0021125|033|nonischemic-frontal impulsivity
C0021125|033|frontotemporal disinhibition
C0021125|033|dementia-related impulsivity
C0021125|033|ad—disinhibition
C0021125|033|ftd—impulsive behavior
C0021125|033|vascular dementia—impulsive
C0021125|033|substance-induced disinhibition
C0021125|033|stimulant-induced impulsivity
C0021125|033|chemo-induced impulsivity
C0021125|033|iatrogenic impulsivity
C0021125|033|ssri-induced impulsivity
C0021125|033|ldopa-induced impulsivity
C0021125|033|pd—impulse control disorder
C0021125|033|pramipexole-induced impulsivity
C0021125|033|dopaminergic impulsivity
C0021125|033|ocd—impulsive symptoms
C0021125|033|borderline impulsivity
C0021125|033|antisocial behavior—impulsivity
C0021125|033|impulsive aggression
C0021125|033|impulsive self-harm
C0021125|033|parasuicidal impulsivity
C0021125|033|sib (self-injurious behavior)
C0021125|033|intermittent explosive episodes
C0021125|033|ied (intermittent explosive disorder)
C0021125|033|dysexecutive impulsivity
C0021125|033|executive function dysregulation
C0021125|033|cognitive impulsivity
C0021125|033|behavioral impulsivity
C0021125|033|motor impulsivity
C0021125|033|verbal impulsivity
C0021125|033|risk-taking behavior
C0021125|033|reckless behavior
C0021125|033|impulsive risk-taking
C0021125|033|failure to inhibit responses
C0021125|033|prepotent response disinhibition
C0021125|033|response inhibition deficit
C0021125|033|dysregulated behavior
C0021125|033|impulse-driven actions
C0021125|033|failure of behavioral restraint
C0021125|033|reward-driven impulsivity
C0021125|033|impulsive motor acts
C0021125|033|short latency responding
C0021125|033|failure to consider consequences
C0021125|033|acting without forethought
C0021125|033|split-second actions
C0021125|033|compromised self-regulation
C0021125|033|poor emotional regulation—impulsivity
C0021125|033|emotion-driven impulsivity
C0021125|033|ir (impulsive responding)
C0021125|033|irb (impulsive/reckless behavior)
C0021125|033|agitated impulsivity
C0021125|033|psychotic impulsivity
C0021125|033|bipolar impulsivity
C0021125|033|schizoaffective—impulsivity
C0021125|033|tic-related impulsivity
C0021125|033|impulsive outbursts
C0021125|033|impulsive speech
C0021125|033|loss of behavioral filter
C0021125|033|uninhibited actions
C0021125|033|loss of frontal lobe inhibition
C0021125|033|impulse dysregulation
C0021125|033|hyperimpulsivity
C0021125|033|pfc dysfunction—impulsivity
C0021125|033|corticobasal syndrome—impulsivity
C0021125|033|impulsive gambling
C0021125|033|compulsive spending—impulsivity
C0021125|033|hypersexuality—impulsivity
C0021125|033|substance binging—impulsivity
C0021125|033|poor delay of gratification
C0021125|033|impaired self-control
C0021125|033|urge-driven behavior
C0021125|033|ictal impulsivity
C0021125|033|seizure-related impulsivity
C0021125|033|irritable impulsivity
C0021125|033|impaired social inhibition
C0021125|033|reckless spending
C0021125|033|rage attacks
C0021125|033|sudden aggressive acts
C0021125|033|reckless driving
C0021125|033|impulsive shoplifting
C0021125|033|pathological impulsivity
C0021125|033|labile impulsivity
C0021125|033|transient disinhibition
C0021125|033|acute-onset disinhibition
C0021125|033|persistent impulsivity
C0021125|033|perseverative impulsivity
C0021125|033|interactive impulsivity
C0021125|033|adolescent impulsivity
C0021125|033|emotional disinhibition
C0021125|033|late-life impulsivity
C0021125|033|childhood impulsivity
C0021125|033|neurocognitive impulsivity
C0021125|033|neurobehavioral disinhibition
C0021125|033|postictal impulsivity
C0021125|033|parkinsonian impulsivity
C0021125|033|impulsive spending
C0021125|033|dysinhibition syndrome
C0021125|033|medication-induced impulsivity
C0021125|033|personality disorder—impulsivity
C0021125|033|impulsive suicidal behavior
C0021125|033|impulsive substance use
C0021125|033|alcohol-related impulsivity
C0021125|033|cns disorder—impulsivity
C0021125|033|chronic impulsivity
C0021125|033|executive system breakdown
C0021125|033|delay aversion
C0021125|033|frontal dysexecutive syndrome
C0021125|033|neurological impulsivity
C0021125|033|psychiatric impulsivity
C0021125|033|primary impulsivity
C0021125|033|secondary impulsivity
C0021125|033|disinhibition (psych/neuro)
C0021125|033|limbic impulsivity
C0021125|033|subcortical impulsivity
C0021125|033|posttraumatic impulsivity
C0021125|033|tbi—impulse control disorder
C0021125|033|impulsive sexual behavior
C0021125|033|shallow decision making
C0021125|033|prefrontal disinhibition
C0021125|033|hyperkinetic impulsivity
C0021125|033|impulsive binge eating
C0021125|033|psychostimulant-induced impulsivity
C0021125|033|parkinsonism—impulsivity
C0021125|033|ftd—behavioral disinhibition
C0021125|033|sud—impulsivity
C0021125|033|emotionally labile—impulsive
C0021125|033|mood-congruent impulsivity
C0021125|033|obsessive-impulsive behavior
C0021125|033|affective impulsivity
C0021125|033|paroxysmal impulsivity
C0021125|033|frontosubcortical impulsivity
C2748208|033|poor executive function
C2748208|033|impaired executive function
C2748208|033|executive dysfunction
C2748208|033|ef deficits
C2748208|033|executive impairment
C2748208|033|deficits in executive function
C2748208|033|executive fx deficits
C2748208|033|executive fx impairment
C2748208|033|dysfunctional executive function
C2748208|033|frontal lobe dysfunction
C2748208|033|frontal executive dysfunction
C2748208|033|executive cognitive deficit
C2748208|033|reduced executive capacity
C2748208|033|impaired ef
C2748208|033|ef impairment
C2748208|033|executive processing deficits
C2748208|033|decreased executive function
C2748208|033|frontal syndrome
C2748208|033|executive skill deficits
C2748208|033|executive control deficit
C2748208|033|impaired cognitive flexibility
C2748208|033|frontally-mediated impairment
C2748208|033|dysexecutive syndrome
C2748208|033|executive system dysfunction
C2748208|033|pfc impairment
C2748208|033|executive performance deficit
C2748208|033|executive control impairment
C2748208|033|cognitive control problems
C2748208|033|loss of executive function
C2748208|033|executive capacity loss
C2748208|033|impaired planning ability
C2748208|033|disorganized thinking
C2748208|033|working memory deficits
C2748208|033|frontal deficits
C2748208|033|frontostriatal dysfunction
C2748208|033|frontosubcortical impairment
C2748208|033|frontal-executive disorder
C2748208|033|frontal executive impairment
C2748208|033|executive fxn problems
C2748208|033|executive dysfunction d/t ad
C2748208|033|executive dysfunction in ftd
C2748208|033|vascular executive dysfunction
C2748208|033|executive dysfunction post-tbi
C2748208|033|executive dysfunction in schizophrenia
C2748208|033|executive dysfunction in mdd
C2748208|033|executive dysfunction in cte
C2748208|033|impaired executive network
C2748208|033|deficient executive processing
C2748208|033|decreased executive skills
C2748208|033|executive attention deficits
C2748208|033|frontal impairment
C2748208|033|executive d/o
C2748208|033|dysexecutive d/o
C2748208|033|frontal lobe syndrome
C2748208|033|impaired task switching
C2748208|033|dysregulated executive function
C2748208|033|impaired ability to plan
C2748208|033|organizing deficits
C2748208|033|sequencing deficits
C2748208|033|inhibition deficit
C2748208|033|problem-solving deficits
C2748208|033|impaired cognitive control
C2748208|033|executive problem
C2748208|033|executive planning difficulties
C2748208|033|loss of executive skills
C2748208|033|frontal circuit impairment
C2748208|033|executive fx difficulty
C2748208|033|executive fxn disruption
C2748208|033|impaired goal-directed behavior
C2748208|033|frontal-subcortical dysfunction
C2748208|033|frontally-based impairment
C2748208|033|pfc d/o
C2748208|033|executive domain impairment
C2748208|033|executive cognitive impairment
C2748208|033|impaired conceptualization
C2748208|033|executive network disruption
C2748208|033|executive impairment w/ vascular etiology
C2748208|033|executive syndrome
C2748208|033|executive control d/o
C2748208|033|abi-related executive dysfunction
C2748208|033|post-stroke executive deficits
C2748208|033|executive dysfunction in svd
C2748208|033|executive impairment secondary to frontal tumor
C2748208|033|executive fxn disorder
C2748208|033|executive processing impairment
C2748208|033|frontal executive deficits
C2748208|033|impaired set-shifting
C2748208|033|executive d/o nos
C2748208|033|executive fxn nos
C2748208|033|impairment in executive abilities
C2748208|033|executive pathway impairment
C2748208|033|dysexecutive pattern
C2748208|033|frontal dysexecutive syndrome
C2748208|033|frontal-executive deficits
C2748208|033|impaired response inhibition
C2748208|033|executive attention impairment
C2748208|033|pfc circuit dysfunction
C2748208|033|cognitive executive dysfunction
C2748208|033|defective executive function
C2748208|033|subcortical executive deficits
C2748208|033|frontal executive domain deficit
C2748208|033|disrupted executive function
C2748208|033|executive dysfunction s/p cva
C2748208|033|executive control failure
C2748208|033|executive dysfunction in adhd
C2748208|033|executive function weaknesses
C2748208|033|executive function disorder
C2748208|033|impaired higher-order control
C2748208|033|executive function abnormality
C2748208|033|executive function underfunction
C2748208|033|executive dysfunction nos
C2748208|033|frontal cognitive impairment
C2748208|033|dysexecutive impairment
C0751295|033|memory loss
C0751295|033|amnestic syndrome
C0751295|033|amnesia
C0751295|033|anterograde amnesia
C0751295|033|retrograde amnesia
C0751295|033|transient global amnesia
C0751295|033|short-term memory loss
C0751295|033|long-term memory loss
C0751295|033|memory impairment
C0751295|033|impaired memory
C0751295|033|cognitive impairment
C0751295|033|cognitive decline
C0751295|033|dementia
C0751295|033|ad
C0751295|033|alzheimer's disease
C0751295|033|vascular dementia
C0751295|033|multi-infarct dementia
C0751295|033|mild cognitive impairment
C0751295|033|mci
C0751295|033|age-associated memory impairment
C0751295|033|post-traumatic amnesia
C0751295|033|traumatic brain injury-related amnesia
C0751295|033|tbi-associated amnesia
C0751295|033|wernicke-korsakoff syndrome
C0751295|033|korsakoff amnesia
C0751295|033|alcohol-related amnesia
C0751295|033|chemo brain
C0751295|033|chemotherapy-induced cognitive impairment
C0751295|033|vascular amnestic syndrome
C0751295|033|hypoxic-ischemic memory loss
C0751295|033|stroke-related memory loss
C0751295|033|postictal amnesia
C0751295|033|epileptic amnesia
C0751295|033|tia-induced memory loss
C0751295|033|tia-related amnesia
C0751295|033|metabolic encephalopathy with memory loss
C0751295|033|encephalopathic memory disturbance
C0751295|033|delirium with impaired recall
C0751295|033|disorientation
C0751295|033|forgetfulness
C0751295|033|poor recall
C0751295|033|poor memory
C0751295|033|difficulty remembering
C0751295|033|loss of memory
C0751295|033|prion disease with memory loss
C0751295|033|creutzfeldt-jakob related memory loss
C0751295|033|frontotemporal dementia with memory deficits
C0751295|033|parkinson's dementia with memory impairment
C0751295|033|lewy body dementia with amnesia
C0751295|033|hiv-associated neurocognitive disorder with memory loss
C0751295|033|ppa with memory involvement
C0751295|033|primary progressive aphasia with memory deficit
C0751295|033|mild amnestic changes
C0751295|033|remote memory loss
C0751295|033|recent memory loss
C0751295|033|febrile amnesia
C0751295|033|post-anoxic amnesia
C0751295|033|toxic encephalopathy with memory loss
C0751295|033|drug-induced amnesia
C0751295|033|medication-related memory loss
C0751295|033|anoxic brain injury-related memory loss
C0751295|033|limbic encephalitis with memory loss
C0751295|033|paraneoplastic limbic encephalitis with amnesia
C0751295|033|autoimmune encephalopathy with memory impairment
C0751295|033|hypoglycemic memory loss
C0751295|033|postictal confusion with amnesia
C0751295|033|infectious encephalopathy with amnesia
C0751295|033|hse memory loss
C0751295|033|herpes simplex encephalitis–related amnesia
C0751295|033|amnestic mild cognitive impairment
C0751295|033|amnestic mci
C0751295|033|global amnesia
C0751295|033|partial amnesia
C0751295|033|focal memory deficit
C0751295|033|subcortical amnesia
C0751295|033|hippocampal amnesia
C0751295|033|amygdalar memory loss
C0751295|033|psychiatric amnesia
C0751295|033|dissociative amnesia
C0751295|033|functional amnesia
C0751295|033|psychogenic amnesia
C0751295|033|hysterical amnesia
C0751295|033|trauma-induced memory loss
C0751295|033|concussion-related amnesia
C0751295|033|blackouts
C0751295|033|confabulatory memory disorder
C0751295|033|confabulation
C0751295|033|mild memory deficit
C0751295|033|significant memory impairment
C0751295|033|progressive memory loss
C0751295|033|chronic memory loss
C0751295|033|paroxysmal amnesia
C0751295|033|acute amnestic episode
C0751295|033|acute memory loss
C0751295|033|episodic memory loss
C0751295|033|semantic memory loss
C0751295|033|working memory deficit
C0751295|033|memory disturbance
C0751295|033|impaired recall
C0751295|033|impaired retention
C0751295|033|defective memory
C0751295|033|failing memory
C0751295|033|loss of retention
C0751295|033|historical amnesia
C0751295|033|anterograde deficit
C0751295|033|retrograde deficit
C0751295|033|ptsd-related amnesia
C0751295|033|stress-induced amnesia
C0751295|033|functional memory loss
C0751295|033|substance-induced memory loss
C0751295|033|prescribed medication-associated amnesia
C0751295|033|amnesia nos
C0751295|033|dementia-related memory loss
C0751295|033|cpm-related memory loss
C0751295|033|central pontine myelinolysis with amnesia
C0751295|033|tumor-related memory loss
C0751295|033|encephalopathic memory defect
C0751295|033|icu-acquired memory deficit
C0751295|033|icu delirium with impaired memory
C0751295|033|nonconvulsive status with amnesia
C0751295|033|nonconvulsive seizure with memory loss
C0751295|033|status epilepticus–related amnesia
C0751295|033|memory deficits
C0751295|033|recall difficulties
C0751295|033|early memory decline
C0751295|033|progressive amnestic disorder
C0751295|033|mild dementia with memory impairment
C0751295|033|mixed dementia with memory loss
C0751295|033|hypertensive encephalopathy with amnesia
C0751295|033|multi-etiology memory loss
C0751295|033|peripartum memory loss
C0751295|033|ppcm with memory impairment
C0751295|033|neurodegenerative memory loss
C0751295|033|amyloid-associated memory decline
C0751295|033|postinfectious memory loss
C0751295|033|hereditary amnesia
C0751295|033|genetic memory impairment
C0751295|033|autosomal dominant amnestic syndrome
C0751295|033|tauopathy with memory loss
C0751295|033|trauma-related memory impairment
C0751295|033|sedative-induced amnesia
C0751295|033|benzodiazepine-related amnesia
C0751295|033|anesthesia-associated amnesia
C0751295|033|anterograde memory deficit
C0751295|033|short-term amnesia
C0751295|033|long-term amnesia
C0751295|033|impaired long-term recall
C0751295|033|memory recall deficit
C0751295|033|subacute memory loss
C0751295|033|transient amnesia
C0751295|033|sudden-onset memory loss
C0751295|033|unexplained amnesia
C0751295|033|idiopathic memory loss
C0751295|033|unspecified amnesia
C0751295|033|attentional amnesia
C0751295|033|tia-induced amnesia
C0751295|033|silent infarct with memory loss
C0751295|033|nonischemic memory loss
C0751295|033|ischemic memory loss
C0751295|033|valvular memory loss
C0751295|033|hypertensive memory loss
C0751295|033|amyloid memory loss
C0751295|033|chemo-induced memory loss
C0751295|033|ppcm-associated memory loss
C0751295|033|tachycardia-induced memory loss
C0751295|033|myocarditis-associated memory loss
C0233794|033|memory impairment
C0233794|033|memory loss
C0233794|033|impaired memory
C0233794|033|amnestic syndrome
C0233794|033|amnesia
C0233794|033|memory dysfunction
C0233794|033|decreased memory
C0233794|033|poor memory
C0233794|033|short-term memory loss
C0233794|033|long-term memory loss
C0233794|033|stm loss
C0233794|033|ltm loss
C0233794|033|anterograde amnesia
C0233794|033|retrograde amnesia
C0233794|033|transient global amnesia
C0233794|033|transient amnesia
C0233794|033|memory deficit
C0233794|033|cognitive impairment
C0233794|033|memory disturbance
C0233794|033|deficit of recall
C0233794|033|recall impairment
C0233794|033|encoding deficit
C0233794|033|retrieval deficit
C0233794|033|executive memory dysfunction
C0233794|033|working memory impairment
C0233794|033|working memory deficit
C0233794|033|impaired recall
C0233794|033|impaired retention
C0233794|033|dementia
C0233794|033|early dementia
C0233794|033|amnestic mci
C0233794|033|mci
C0233794|033|mild cognitive impairment
C0233794|033|vuci (vascular unrelated cognitive impairment)
C0233794|033|vci (vascular cognitive impairment)
C0233794|033|post-stroke memory loss
C0233794|033|ischemic memory loss
C0233794|033|vascular memory deficit
C0233794|033|nonischemic memory loss
C0233794|033|hypoxic memory impairment
C0233794|033|hypoxic brain injury with memory loss
C0233794|033|postencephalitic memory loss
C0233794|033|encephalopathic memory deficit
C0233794|033|tbi memory loss
C0233794|033|post-concussive amnesia
C0233794|033|concussion-related memory loss
C0233794|033|chemotherapy-induced memory impairment
C0233794|033|chemo brain
C0233794|033|radiation-induced memory deficit
C0233794|033|alcohol-related memory impairment
C0233794|033|wernicke-korsakoff amnesia
C0233794|033|thiamine deficiency–related memory loss
C0233794|033|alzheimer's-related memory loss
C0233794|033|ad-associated memory loss
C0233794|033|ftd memory loss
C0233794|033|frontotemporal dementia memory deficit
C0233794|033|pca memory impairment
C0233794|033|posterior cortical atrophy with memory loss
C0233794|033|lewy body dementia–associated memory loss
C0233794|033|lbd memory loss
C0233794|033|parkinson's with memory impairment
C0233794|033|pd memory deficit
C0233794|033|multiple sclerosis with memory loss
C0233794|033|ms-related memory impairment
C0233794|033|huntington’s chorea with memory loss
C0233794|033|amyloid-related memory impairment
C0233794|033|neurodegenerative memory loss
C0233794|033|iatrogenic memory deficit
C0233794|033|medication-related memory loss
C0233794|033|benzo-induced memory loss
C0233794|033|steroid-induced cognitive impairment
C0233794|033|psychiatric memory loss
C0233794|033|ptsd-related memory gap
C0233794|033|depressive pseudodementia
C0233794|033|anxiety-related memory impairment
C0233794|033|stress-induced memory deficit
C0233794|033|age-associated memory impairment
C0233794|033|presbycognitive change
C0233794|033|elderly memory decline
C0233794|033|mild memory decline
C0233794|033|subjective memory complaint
C0233794|033|forgetfulness
C0233794|033|recent memory deficit
C0233794|033|remote memory deficit
C0233794|033|remote memory impairment
C0233794|033|recognition impairment
C0233794|033|impaired knowledge retention
C0233794|033|deficient recall
C0233794|033|blackout (memory)
C0233794|033|global amnesia
C0233794|033|functional amnesia
C0233794|033|psychogenic amnesia
C0233794|033|dissociative amnesia
C0233794|033|hysterical amnesia
C0233794|033|traumatic amnesia
C0233794|033|reversible memory impairment
C0233794|033|irreversible memory impairment
C0233794|033|progressive memory loss
C0233794|033|episodic memory loss
C0233794|033|semantic memory loss
C0233794|033|immediate memory deficit
C0233794|033|delayed recall loss
C0233794|033|impaired new learning
C0233794|033|learning disability (acquired)
C0233794|033|impaired memory acquisition
C0233794|033|anterograde deficit
C0233794|033|retrograde deficit
C0233794|033|amnesic syndrome
C0233794|033|drug-induced amnesia
C0233794|033|toxic encephalopathy with memory loss
C0233794|033|metabolic encephalopathy with memory impairment
C0233794|033|autoimmune encephalitis–associated memory loss
C0233794|033|limbic encephalitis–associated memory loss
C0233794|033|temporal lobe memory deficit
C0233794|033|frontal lobe memory deficit
C0233794|033|medial temporal amnesia
C0233794|033|devastating memory loss
C0233794|033|attentional memory deficit
C0233794|033|ppcm-related cognitive deficit
C0233794|033|post-infectious cognitive impairment
C0233794|033|covid-related cognitive impairment
C0233794|033|long covid memory issues
C0233794|033|hiv-associated neurocognitive memory loss
C0233794|033|cjd memory loss
C0233794|033|prion-related memory deficit
C0233794|033|chronic memory loss
C0233794|033|acute memory loss
C0233794|033|subacute memory loss
C0233794|033|abrupt memory deficit
C0233794|033|persistent memory impairment
C0233794|033|fluctuating memory impairment
C0233794|033|paraneoplastic-related memory deficit
C0233794|033|seizure-associated amnesia
C0233794|033|postictal amnesia
C0233794|033|postictal confusion with memory loss
C0233794|033|epileptic amnesia
C0233794|033|epilepsy-related memory impairment
C0233794|033|temporal lobe epilepsy amnesia
C0233794|033|tle-associated memory loss
C0233794|033|atrial fibrillation–related memory loss
C0233794|033|af-related cognitive deficit
C0233794|033|hypertensive memory deficit
C0233794|033|cardiac memory loss
C0233794|033|chf-related memory impairment
C0233794|033|heart failure–associated cognitive impairment
C0233794|033|tachycardia-induced cognitive dysfunction
C0233794|033|tci-related memory loss
C0233794|033|neuropathic memory deficit
C0233794|033|cortical memory impairment
C0233794|033|subcortical memory impairment
C0233794|033|hie-related memory loss
C0233794|033|hypoxic-ischemic encephalopathy with memory loss
C0233794|033|hypoperfusion-related cognitive deficit
C0233794|033|dialysis dementia
C0233794|033|renal failure-related memory loss
C0233794|033|hepatic encephalopathy with memory deficit
C0233794|033|liver failure–related cognitive disorder
C0233794|033|systemic illness–related memory impairment
C0233794|033|delirium-associated amnesia
C0233794|033|icu-related memory deficit
C0233794|033|post-surgical memory loss
C0233794|033|perioperative amnesia
C0233794|033|critical illness–associated cognitive impairment
C0233407|033|disoriented
C0233407|033|disorientation
C0233407|033|ams
C0233407|033|altered mental status
C0233407|033|confusion
C0233407|033|confused
C0233407|033|delirium
C0233407|033|delirious
C0233407|033|mental status changes
C0233407|033|acute confusional state
C0233407|033|waxing and waning mental status
C0233407|033|disorganized thought process
C0233407|033|disorganized thought
C0233407|033|incoherent
C0233407|033|encephalopathy
C0233407|033|acute encephalopathy
C0233407|033|lethargy
C0233407|033|obtunded
C0233407|033|clouded sensorium
C0233407|033|mental clouding
C0233407|033|senile confusion
C0233407|033|acute mental status change
C0233407|033|altered level of consciousness
C0233407|033|near-syncope with confusion
C0233407|033|post-ictal confusion
C0233407|033|toxic-metabolic encephalopathy
C0233407|033|confusional state
C0233407|033|transient confusion
C0233407|033|acute organic brain syndrome
C0233407|033|disorientation to time
C0233407|033|disorientation to place
C0233407|033|disorientation to person
C0233407|033|chrono-disorientation
C0233407|033|spatial disorientation
C0233407|033|person-place-time disorientation
C0233407|033|aox1
C0233407|033|aox2
C0233407|033|not aox3
C0233407|033|not alert and oriented
C0233407|033|poor orientation
C0233407|033|oriented x1
C0233407|033|oriented x2
C0233407|033|oriented x0
C0233407|033|diminished awareness
C0233407|033|no orientation
C0233407|033|stuporous
C0233407|033|disoriented behavior
C0233407|033|mental fog
C0233407|033|altered sensorium
C0233407|033|disoriented to surroundings
C0233407|033|cognitive dysfunction
C0233407|033|cognitive impairment
C0233407|033|acute mental confusion
C0233407|033|waxing/waning orientation
C0233407|033|episodes of confusion
C0233407|033|vague mentation
C0233407|033|inattentive
C0233407|033|memory lapse with confusion
C0233407|033|icu delirium
C0233407|033|hosp. delirium
C0233407|033|sun-downing
C0233407|033|sundowning
C0233407|033|critical illness encephalopathy
C0233407|033|hepatic encephalopathy
C0233407|033|uremic encephalopathy
C0233407|033|metabolic encephalopathy
C0233407|033|hypoxic encephalopathy
C0233407|033|septic encephalopathy
C0233407|033|postictal state
C0233407|033|confusional episode
C0233407|033|transient disorientation
C0233407|033|altered awareness
C0233407|033|impaired orientation
C0233407|033|o/e: disoriented
C0233407|033|aox1 (person)
C0233407|033|aox1 (place)
C0233407|033|aox1 (time)
C0233407|033|unoriented
C0233407|033|not oriented
C0233407|033|losing orientation
C0233407|033|fluctuating mental status
C0233407|033|acute onset confusion
C0233407|033|dementia-related confusion
C0233407|033|psychotic disorganization
C0233407|033|mental status waxing/waning
C0233407|033|short-term confusion
C0233407|033|periodic confusion
C0233407|033|post-operative confusion
C0233407|033|icu psychosis
C0233407|033|post-op delirium
C0233407|033|chemotherapy-induced delirium
C0233407|033|drug-induced confusion
C0233407|033|intoxication delirium
C0233407|033|withdrawal-related confusion
C0233407|033|alcoholic encephalopathy
C0233407|033|wernicke's encephalopathy
C0233407|033|delirium tremens
C0233407|033|tachycardia-induced confusion
C0233407|033|sepsis-induced ams
C0233407|033|infection-related altered mentation
C0233407|033|ppcm-related ams
C0233407|033|myocarditis delirium
C0233407|033|ischemic encephalopathy
C0233407|033|stroke-related confusion
C0233407|033|tia-related ams
C0233407|033|vascular dementia w/ confusion
C0233407|033|valvular disease ams
C0233407|033|hypertensive encephalopathy
C0233407|033|amyloid encephalopathy
C0233407|033|hypoglycemia with confusion
C0233407|033|hyperglycemic confusion
C0233407|033|dka-related ams
C0233407|033|hhs with disorientation
C0233407|033|hypercapnic encephalopathy
C0233407|033|co2 narcosis
C0233407|033|hypoxemic confusion
C0233407|033|anoxic encephalopathy
C0233407|033|thiamine-deficiency encephalopathy
C0233407|033|nonconvulsive status ams
C0233407|033|paraneoplastic encephalopathy
C0233407|033|tumor-related confusion
C0233407|033|brain metastasis ams
C0233407|033|space-occupying lesion ams
C0233407|033|subdural hematoma with confusion
C0233407|033|sah with disorientation
C0233407|033|traumatic brain injury ams
C0233407|033|mild cognitive impairment with confusion
C0233407|033|multifactorial ams
C0233407|033|confusional syndrome
C0233407|033|encephalopathic state
C0233407|033|organic brain syndrome
C0233407|033|momentary confusion
C0233407|033|low arousal state
C0233407|033|poor mentation
C0233407|033|encephalopathic changes
C0233407|033|delayed mentation
C0233407|033|nonresponsive with confusion
C0233407|033|unresponsive with confusion
C0233407|033|somnolent
C0233407|033|stupor with disorientation
C0233407|033|not alert
C0233407|033|disorganized mentation
C0233407|033|psychomotor disorientation
C0233407|033|cerebral dysfunction
C0233407|033|disoriented to environment
C0233407|033|no orientation to date
C0233407|033|no orientation to location
C0233407|033|acute confusion state
C0233407|033|hyperactive delirium
C0233407|033|hypoactive delirium
C0233407|033|mixed delirium
C0233407|033|fluctuating orientation
C0233407|033|confused on exam
C0233407|033|disoriented on assessment
C0233407|033|not oriented on exam
C0233407|033|o/e: confused
C0233407|033|patient confused
C0233407|033|pt confused
C0233407|033|pt disoriented
C0233407|033|aox0
C0233407|033|unaware of time/place
C0233407|033|disorientation to situation
C0233407|033|not oriented to time
C0233407|033|not oriented to place
C0233407|033|not oriented to self
C0233407|033|not oriented to situation
C0233407|033|orientation deficit
C0233407|033|impaired consciousness
C0233407|033|poor cognition
C0233407|033|acute altered consciousness
C0233407|033|mental slowing
C0233407|033|ams of unclear etiology
C0233407|033|global confusion
C0233407|033|cerebral confusion
C0233407|033|organic confusion
C0233407|033|cns dysfunction with confusion
C0233407|033|mental status alteration
C0233407|033|loss of orientation
C0233407|033|labile orientation
C0233407|033|impaired mentation
C0233407|033|not ao
C0233407|033|disturbed consciousness
C0015676|033|mental fatigue
C0015676|033|cognitive fatigue
C0015676|033|cognitive exhaustion
C0015676|033|cognitive weariness
C0015676|033|psychic fatigue
C0015676|033|psychic exhaustion
C0015676|033|psychic weariness
C0015676|033|neurofatigue
C0015676|033|neurocognitive fatigue
C0015676|033|mental exhaustion
C0015676|033|mental weariness
C0015676|033|mental tiredness
C0015676|033|cognitive tiredness
C0015676|033|psychological fatigue
C0015676|033|brain fatigue
C0015676|033|brain fog
C0015676|033|brain tiredness
C0015676|033|mental sluggishness
C0015676|033|decreased mental stamina
C0015676|033|neural fatigue
C0015676|033|cognitive slowing
C0015676|033|decreased cognitive endurance
C0015676|033|decreased concentration endurance
C0015676|033|loss of mental stamina
C0015676|033|reduced cognitive capacity
C0015676|033|subjective cognitive fatigue
C0015676|033|cerebral fatigue
C0015676|033|cortical fatigue
C0015676|033|chemo brain
C0015676|033|chemo-induced cognitive fatigue
C0015676|033|chemo-related brain fog
C0015676|033|crf (cancer-related fatigue)
C0015676|033|crcf (cancer-related cognitive fatigue)
C0015676|033|ms-related cognitive fatigue
C0015676|033|stroke-related mental fatigue
C0015676|033|ischemic cognitive fatigue
C0015676|033|nonischemic mental fatigue
C0015676|033|tbi-related mental fatigue
C0015676|033|postconcussive fatigue
C0015676|033|neurological fatigue
C0015676|033|als-related cognitive fatigue
C0015676|033|pd-related cognitive fatigue
C0015676|033|dementia-related fatigue
C0015676|033|depression-related fatigue
C0015676|033|post-stroke cognitive fatigue
C0015676|033|cfs-related mental fatigue
C0015676|033|chronic fatigue syndrome mental exhaustion
C0015676|033|primary fatigue of ms
C0015676|033|encephalopathic fatigue
C0015676|033|paraneoplastic fatigue
C0015676|033|autoimmune encephalitis cognitive fatigue
C0015676|033|ra-related mental fatigue
C0015676|033|lupus-related cognitive fatigue
C0015676|033|post-viral fatigue
C0015676|033|long covid brain fog
C0015676|033|pasc cognitive fatigue
C0015676|033|mental lassitude
C0015676|033|mental depletion
C0015676|033|attention fatigue
C0015676|033|executive fatigue
C0015676|033|decision fatigue
C0015676|033|sustained attention impairment
C0015676|033|mental stamina loss
C0015676|033|cognitive burnout
C0015676|033|mental burnout
C0015676|033|neuropsychiatric fatigue
C0015676|033|postictal fatigue
C0015676|033|post-seizure cognitive fatigue
C0015676|033|fibro fog
C0015676|033|fibromyalgia-related cognitive fatigue
C0015676|033|psychiatric fatigue
C0015676|033|schizophrenia-related cognitive fatigue
C0015676|033|bipolar-related cognitive fatigue
C0015676|033|ptsd-related cognitive fatigue
C0015676|033|csf (chronic symptom fatigue)
C0015676|033|chronic illness fatigue
C0015676|033|pots-related cognitive fatigue
C0015676|033|orthostatic cognitive fatigue
C0015676|033|dysautonomia fatigue
C0015676|033|anemia-related mental fatigue
C0015676|033|metabolic fatigue
C0015676|033|liver disease-related mental fatigue
C0015676|033|ckd-related cognitive fatigue
C0015676|033|dialysis-related cognitive fatigue
C0015676|033|hypothyroidism-related cognitive fatigue
C0015676|033|sle mental fatigue
C0015676|033|immune-mediated cognitive fatigue
C0015676|033|cancer brain fog
C0015676|033|brain fatigue syndrome
C0015676|033|postviral fatigue syndrome
C0015676|033|vaccination-related cognitive fatigue
C0015676|033|viral encephalitis-related fatigue
C0015676|033|substance-induced mental fatigue
C0015676|033|medication-induced cognitive fatigue
C0015676|033|drug-induced cognitive fatigue
C0015676|033|cognitive malaise
C0015676|033|nonrestorative cognitive fatigue
C0015676|033|fatigued cognition
C0015676|033|overtired mental state
C0015676|033|prolonged cognitive fatigue
C0015676|033|prolonged mental exhaustion
C0015676|033|work-related mental fatigue
C0015676|033|post-work mental exhaustion
C0015676|033|shift work-related mental fatigue
C0015676|033|vhf (viral hemorrhagic fever) related fatigue
C0015676|033|covid-19 related brain fog
C0015676|033|fatigue of central origin
C0015676|033|central fatigue
C0015676|033|pervasive cognitive fatigue
C0015676|033|psychomotor slowing
C0015676|033|cognitive inefficiency
C0015676|033|mental inefficiency
C0015676|033|cognitive drain
C0015676|033|mental drain
C0015676|033|cognitive depletion
C0015676|033|ptf (post-traumatic fatigue)
C0015676|033|fatigue nos
C0015676|033|subjective mental fatigue
C0015676|033|subjective brain fog
C0015676|033|reduced cognitive throughput
C0015676|033|cognitive wearout
C0015676|033|cognitive clouding
C0015676|033|mental fog
C0015676|033|decreased processing speed
C0015676|033|information processing fatigue
C0015676|033|executive function fatigue
C0015676|033|mental lethargy
C0015676|033|cognitive lethargy
C0015676|033|mental clouding
C0015676|033|cognitive cloudiness
C0015676|033|brain exhaustion
C0015676|033|mental enervation
C0015676|033|cognitive enervation
C0015676|033|loss of mental acuity
C0015676|033|decreased alertness
C0015676|033|sustained attention fatigue
C0015676|033|prolonged attentional fatigue
C0015676|033|prolonged vigilance fatigue
C0015676|033|vigilance decrement
C0015676|033|alertness decline
C0015676|033|delayed mental response
C0015676|033|mental processing delay
C0015676|033|cortical exhaustion
C0015676|033|frontal fatigue
C0015676|033|frontosubcortical fatigue
C0015676|033|psychogenic fatigue
C0015676|033|psychological exhaustion
C0015676|033|psychological tiredness
C0015676|033|occupational cognitive fatigue
C0015676|033|occupational brain fatigue
C0015676|033|task-related mental fatigue
C0015676|033|task-induced fatigue
C0015676|033|workload-related cognitive fatigue
C0015676|033|shiftwork fatigue
C0015676|033|driver fatigue (mental)
C0015676|033|operator mental fatigue
C0015676|033|performance fatigue
C0015676|033|mental overexertion
C0015676|033|cerebral exhaustion
C0015676|033|cognitive slowing syndrome
C0015676|033|effort fatigue
C0015676|033|expended cognitive reserves
C0015676|033|decreased cognitive reserves
C0015676|033|mental performance decrement
C0015676|033|mental function decrement
C0015676|033|ppcs-related fatigue
C0015676|033|post-tia cognitive fatigue
C0015676|033|hiv-associated neurocognitive fatigue
C0015676|033|aids-related cognitive fatigue
C0015676|033|immunotherapy-related brain fog
C0015676|033|antiviral-induced cognitive fatigue
C0015676|033|anticholinergic-related cognitive fatigue
C0015676|033|steroid-related cognitive fatigue
C0015676|033|anti-epileptic-induced cognitive fatigue
C0015676|033|antipsychotic-related cognitive fatigue
C0015676|033|depressogenic fatigue
C0015676|033|icu-related cognitive fatigue
C0015676|033|post-icu fatigue
C0015676|033|post-hospitalization mental fatigue
C0015676|033|sleep deprivation-related mental fatigue
C0015676|033|insomnia-related cognitive fatigue
C0015676|033|sleep disorder mental fatigue
C0015676|033|hypersomnia mental fatigue
C0015676|033|shiftwork disorder-related mental fatigue
C0015676|033|disrupted circadian cognitive fatigue
C0015676|033|nocturnal cognitive fatigue
C0015676|033|daytime cognitive fatigue
C0029227|033|delirium
C0029227|033|acute confusional state
C0029227|033|acute brain syndrome
C0029227|033|acute encephalopathy
C0029227|033|icu psychosis
C0029227|033|toxic encephalopathy
C0029227|033|substance-induced delirium
C0029227|033|alcohol withdrawal delirium
C0029227|033|delirium tremens
C0029227|033|hyperactive delirium
C0029227|033|hypoactive delirium
C0029227|033|mixed delirium
C0029227|033|dementia
C0029227|033|major neurocognitive disorder
C0029227|033|minor neurocognitive disorder
C0029227|033|neurocognitive disorder nos
C0029227|033|primary degenerative dementia
C0029227|033|senile dementia
C0029227|033|presenile dementia
C0029227|033|senile cortical degeneration
C0029227|033|multi-infarct dementia
C0029227|033|vascular dementia
C0029227|033|ischemic vascular dementia
C0029227|033|nonischemic dementia
C0029227|033|subcortical dementia
C0029227|033|frontotemporal dementia
C0029227|033|pick's disease
C0029227|033|lewy body dementia
C0029227|033|parkinson’s disease dementia
C0029227|033|alzheimer’s disease
C0029227|033|ad
C0029227|033|alzheimers type dementia
C0029227|033|dementia with behavioral disturbance
C0029227|033|dementia with psychosis
C0029227|033|dementia with delusions
C0029227|033|dementia with agitation
C0029227|033|dementia with depression
C0029227|033|aids dementia complex
C0029227|033|hiv-associated dementia
C0029227|033|chemo-induced cognitive impairment
C0029227|033|chemotherapy-related cognitive dysfunction
C0029227|033|chemo brain
C0029227|033|alcohol-related dementia
C0029227|033|wernicke-korsakoff syndrome
C0029227|033|korsakoff dementia
C0029227|033|wernicke’s encephalopathy
C0029227|033|normal pressure hydrocephalus
C0029227|033|nph
C0029227|033|post-stroke dementia
C0029227|033|postinfectious dementia
C0029227|033|pandas encephalopathy
C0029227|033|creutzfeldt-jakob disease
C0029227|033|prion disease dementia
C0029227|033|huntington’s disease dementia
C0029227|033|hd dementia
C0029227|033|rapidly progressive dementia
C0029227|033|progressive supranuclear palsy dementia
C0029227|033|depression-related cognitive impairment
C0029227|033|pseudo-dementia
C0029227|033|amnestic disorder
C0029227|033|amnestic syndrome
C0029227|033|amnestic mci
C0029227|033|anoxic brain injury dementia
C0029227|033|hypoxic-ischemic encephalopathy
C0029227|033|down syndrome dementia
C0029227|033|ds dementia
C0029227|033|mild cognitive impairment
C0029227|033|mci
C0029227|033|age-related cognitive decline
C0029227|033|cognitive disorder nos
C0029227|033|organic brain syndrome
C0029227|033|organic mental disorder
C0029227|033|cognitive dysfunction
C0029227|033|cognitive decline
C0029227|033|chronic confusional state
C0029227|033|global cognitive impairment
C0029227|033|memory loss
C0029227|033|short-term memory loss
C0029227|033|long-term memory loss
C0029227|033|executive dysfunction
C0029227|033|aphasic dementia
C0029227|033|primary progressive aphasia
C0029227|033|semantic dementia
C0029227|033|logopenic progressive aphasia
C0029227|033|agrammatic aphasia
C0029227|033|cadasil dementia
C0029227|033|amyloid angiopathy-related dementia
C0029227|033|posterior cortical atrophy
C0029227|033|binswanger's disease
C0029227|033|thalamic dementia
C0029227|033|corticobasal degeneration dementia
C0029227|033|cbd dementia
C0029227|033|marchiafava-bignami disease
C0029227|033|menstrual-related cognitive changes
C0029227|033|steroid-induced cognitive dysfunction
C0029227|033|medication-induced encephalopathy
C0029227|033|paraneoplastic encephalopathy
C0029227|033|autoimmune encephalopathy
C0029227|033|anti-nmda receptor encephalitis
C0029227|033|syphilitic dementia
C0029227|033|neurosyphilis dementia
C0029227|033|wilson’s disease dementia
C0029227|033|copper-related cognitive disorder
C0029227|033|b12 deficiency dementia
C0029227|033|hypothyroid dementia
C0029227|033|hypoglycemic encephalopathy
C0029227|033|hypoparathyroidism cognitive dysfunction
C0029227|033|hypercalcemia cognitive impairment
C0029227|033|postictal confusion
C0029227|033|chronic traumatic encephalopathy
C0029227|033|ptsd-related cognitive disorder
C0029227|033|cognitive impairment nos
C0029227|033|transient global amnesia
C0029227|033|fahr's syndrome dementia
C0029227|033|basal ganglia dementia
C0029227|033|epileptic encephalopathy
C0029227|033|retrospective amnesia
C0029227|033|anterograde amnesia
C0029227|033|retrograde amnesia
C0029227|033|secondary dementia
C0029227|033|delirious mania
C0029227|033|steroid psychosis
C0029227|033|icu delirium
C0029227|033|withdrawal delirium
C0029227|033|metabolic encephalopathy
C0029227|033|hepatic encephalopathy
C0029227|033|uremic encephalopathy
C0029227|033|dialysis dementia
C0029227|033|dialysis encephalopathy
C0029227|033|hypoxic encephalopathy
C0029227|033|hypoxic-ischemic brain injury
C0029227|033|acute memory loss
C0029227|033|psychosis with cognitive decline
C0029227|033|behavioral variant dementia
C0029227|033|semantic variant primary progressive aphasia
C0029227|033|nonfluent variant primary progressive aphasia
C0029227|033|progressive nonfluent aphasia
C0029227|033|alzheimer-type psychosis
C0029227|033|mild ncd
C0029227|033|major ncd
C0029227|033|cognitive disorder due to trauma
C0029227|033|postconcussive syndrome cognitive deficit
C0029227|033|residual cognitive deficits
C0029227|033|ppcm cognitive disorder
C0029227|033|postpartum cognitive impairment
C0029227|033|peripartum cognitive disorder
C0029227|033|tachycardia-induced encephalopathy
C0029227|033|valvular-related dementia
C0029227|033|amyloid-related cognitive impairment
C0029227|033|toxic-metabolic encephalopathy
C0029227|033|dementia nos
C0029227|033|senile ncd
C0029227|033|mixed ncd
C0029227|033|age-associated memory impairment
C0029227|033|cortical dementia
C0029227|033|subcortical cognitive disorder
C0029227|033|ischemic encephalopathy
C0029227|033|hypertensive encephalopathy
C0029227|033|cadasil cognitive impairment
C0029227|033|binswanger type ncd
C0029227|033|cerebral amyloid angiopathy cognitive dysfunction
C0009676|033|confusion
C0009676|033|confused
C0009676|033|ams
C0009676|033|altered mental status
C0009676|033|acute confusion
C0009676|033|delirium
C0009676|033|encephalopathy
C0009676|033|acute encephalopathy
C0009676|033|subacute confusion
C0009676|033|disoriented
C0009676|033|disorientation
C0009676|033|impaired consciousness
C0009676|033|clouded sensorium
C0009676|033|impaired awareness
C0009676|033|decreased alertness
C0009676|033|impaired mentation
C0009676|033|drowsy
C0009676|033|obtunded
C0009676|033|lethargic
C0009676|033|waxing/waning level of consciousness
C0009676|033|inattentive
C0009676|033|difficulty following commands
C0009676|033|mental status change
C0009676|033|acute mental status change
C0009676|033|cognitive dysfunction
C0009676|033|cognitive disturbance
C0009676|033|delirious
C0009676|033|somnolent
C0009676|033|fluctuating mental status
C0009676|033|with confusion
C0009676|033|episodes of confusion
C0009676|033|disorganized thinking
C0009676|033|impaired thought process
C0009676|033|slowed thought process
C0009676|033|slowed cognition
C0009676|033|stuporous
C0009676|033|coma
C0009676|033|minimally responsive
C0009676|033|encephalopathic
C0009676|033|toxic/metabolic encephalopathy
C0009676|033|hepatic encephalopathy
C0009676|033|septic encephalopathy
C0009676|033|postictal confusion
C0009676|033|icu delirium
C0009676|033|hypoxic encephalopathy
C0009676|033|wernicke’s encephalopathy
C0009676|033|ischemic encephalopathy
C0009676|033|hypoperfusion encephalopathy
C0009676|033|agitated confusion
C0009676|033|restless and confused
C0009676|033|dementia with acute change
C0009676|033|delirium superimposed on dementia
C0009676|033|waxing/waning cognition
C0009676|033|transient confusion
C0009676|033|acute confusional state
C0009676|033|acd (acute confusional disorder)
C0009676|033|delirium nos
C0009676|033|confusional syndrome
C0009676|033|mixed hypoactive/hyperactive delirium
C0009676|033|perplexed
C0009676|033|pocd (postoperative cognitive dysfunction)
C0009676|033|encephalopathic state
C0009676|033|confusional episode
C0009676|033|psycho-organic syndrome
C0009676|033|cognitive impairment
C0009676|033|delirious state
C0009676|033|decreased cognition
C0009676|033|mental confusion
C0009676|033|acute brain dysfunction
C0009676|033|neurocognitive dysfunction
C0009676|033|incoherent
C0009676|033|psychosis (if used for acute confusion)
C0009676|033|muddled
C0009676|033|muddled thinking
C0009676|033|acute brain failure
C0009676|033|disorganized speech
C0009676|033|delayed response
C0009676|033|impaired attention
C0009676|033|short-term memory loss
C0009676|033|unresponsive (when r/t confusion)
C0009676|033|impaired memory and orientation
C0009676|033|reduced arousal
C0009676|033|fluctuating alertness
C0009676|033|depressed level of consciousness
C0009676|033|hyperactive delirium
C0009676|033|hypoactive delirium
C0009676|033|confusional psychosis
C0009676|033|delirium tremens
C0009676|033|delirium due to substance
C0009676|033|withdrawal delirium
C0009676|033|drug-induced confusion
C0009676|033|chemo-induced confusion
C0009676|033|post-stroke confusion
C0009676|033|tia-related confusion
C0009676|033|incoherent mental status
C0009676|033|spoken incoherence
C0009676|033|mistakes place and time
C0009676|033|impaired executive function
C0009676|033|disordered consciousness
C0009676|033|acute brain syndrome
C0009676|033|transient global amnesia (if confused)
C0009676|033|cns dysfunction
C0009676|033|metabolic confusion
C0009676|033|senile confusion
C0009676|033|delirium due to uti
C0009676|033|hospital-acquired delirium
C0009676|033|pod (postoperative delirium)
C0009676|033|encephalopathy nos
C0009676|033|septic confusion
C0009676|033|disorganized behavior
C0009676|033|acute cognitive impairment
C0009676|033|chronic confusion
C0009676|033|substance-induced confusion
C0009676|033|fluctuating cognition
C0009676|033|distractible
C0009676|033|frontal syndrome
C0009676|033|sundowning
C0009676|033|decreased responsiveness
C0009676|033|confusional state nos
C0009676|033|agitated delirium
C0009676|033|restless mental status
C0009676|033|delirium secondary to infection
C0009676|033|delirium of metabolic origin
C0009676|033|delirium due to hypoxia
C0009676|033|paranoia with confusion
C0009676|033|encephalopathic confusion
C0009676|033|mistakes relatives
C0009676|033|word salad
C0009676|033|rambling speech
C0009676|033|unorganized thought process
C0009676|033|thought disorder
C0009676|033|reduced mentation
C0009676|033|abnormal mentation
C0009676|033|periods of unresponsiveness
C0009676|033|clouding of consciousness
C0009676|033|icu psychosis
C0009676|033|acute organic brain syndrome
C0009676|033|toxic psychosis
C0009676|033|organic psychosis
C0009676|033|paranoid confusion
C0009676|033|impaired judgement
C0009676|033|bilious confusion (rare)
C0009676|033|delayed recall
C0009676|033|memory lapses
C0009676|033|impaired cognitive status
C0009676|033|disoriented to time
C0009676|033|disoriented to place
C0009676|033|disoriented to person
C0009676|033|delays in thought
C0009676|033|thought blocking
C0009676|033|forgetful
C0009676|033|attention deficit
C0009676|033|unusual behavior
C0009676|033|disinhibited
C0009676|033|wandering
C0009676|033|not oriented
C0009676|033|not following commands
C0009676|033|memory disturbance
C0009676|033|confabulating
C0009676|033|semantic paraphasia
C0009676|033|aphasic confusion
C0009676|033|acute on chronic confusion
C0009676|033|episodic confusion
C0009676|033|impaired recall
C0009676|033|executive dysfunction
C0009676|033|new cognitive deficit
C0009676|033|fluency disturbance
C0009676|033|paraphasic errors
C0009676|033|confusional arousal
C0009676|033|psychomotor agitation
C0009676|033|psychomotor retardation
C0009676|033|frontal release signs
C0009676|033|amnesia with confusion
C0009676|033|postictal state
C0009676|033|post-ictal confusion
C0009676|033|acute delirium
C0009676|033|dementia with acute confusion
C0009676|033|loc fluctuation
C0009676|033|fluctuating loc
C0009676|033|perseveration (if confused)
C0009676|033|incoherence
C0009676|033|speech disorganization
C0009676|033|language disturbance
C0009676|033|labile mood (if confused)
C0009676|033|inappropriate affect with confusion
C0009676|033|paraphasic confusion
C0009676|033|organically based confusion
C0009676|033|toxic confusion
C0009676|033|leukoencephalopathic confusion
C0009676|033|drug-related encephalopathy
C0009676|033|viral encephalopathy with confusion
C0009676|033|postoperative confusion
C0009676|033|post-anesthesia confusion
C0009676|033|pse (portosystemic encephalopathy)
C0233414|033|impaired attention
C0233414|033|inattentiveness
C0233414|033|poor attention
C0233414|033|decreased attention
C0233414|033|attention deficit
C0233414|033|attention disturbance
C0233414|033|deficit in attention
C0233414|033|distractibility
C0233414|033|difficulty focusing
C0233414|033|shortened attention span
C0233414|033|distraction
C0233414|033|problems concentrating
C0233414|033|concentration deficit
C0233414|033|impaired concentration
C0233414|033|reduced concentration
C0233414|033|decreased concentration
C0233414|033|difficulty concentrating
C0233414|033|unable to concentrate
C0233414|033|concentration disturbance
C0233414|033|attentional impairment
C0233414|033|fluctuating attention
C0233414|033|labile attention
C0233414|033|poor focus
C0233414|033|impaired focus
C0233414|033|easily distracted
C0233414|033|ad
C0233414|033|inability to sustain attention
C0233414|033|inattention
C0233414|033|selective inattention
C0233414|033|failing to attend
C0233414|033|loc impairment (level of consciousness)
C0233414|033|clouded attention
C0233414|033|clouded consciousness
C0233414|033|diffuse attentional disturbance
C0233414|033|nonpersistent attention
C0233414|033|transient attention loss
C0233414|033|brief attention span
C0233414|033|inattentive state
C0233414|033|wandering attention
C0233414|033|unstable attention
C0233414|033|transient inattention
C0233414|033|attention span impairment
C0233414|033|mental inattentiveness
C0233414|033|failure to focus
C0233414|033|short attention span
C0233414|033|distractible
C0233414|033|attentional deficit
C0233414|033|delirium (if used to mean attention disturbance)
C0233414|033|delirious (as shorthand)
C0233414|033|delirium syndrome
C0233414|033|fluctuating awareness
C0233414|033|hypoactive attention
C0233414|033|aao ×3 poor
C0233414|033|impaired vigilance
C0233414|033|reduced vigilance
C0233414|033|dysexecutive syndrome
C0233414|033|executive dysfunction
C0233414|033|non-focal attentional deficit
C0233414|033|subcortical attention impairment
C0233414|033|ischemic attention disturbance
C0233414|033|metabolic attention impairment
C0233414|033|hepatic attention disturbance
C0233414|033|toxic attention impairment
C0233414|033|infectious attention deficit
C0233414|033|delirium d/t infection
C0233414|033|delirium d/t uti
C0233414|033|delirium d/t sepsis
C0233414|033|chemo-induced attention deficit
C0233414|033|attention deficit secondary to tbi
C0233414|033|encephalopathic attention deficit
C0233414|033|drug-induced inattention
C0233414|033|alcohol-related inattention
C0233414|033|paraneoplastic attention deficit
C0233414|033|cancer-related attention deficit
C0233414|033|neurologic attention deficit
C0233414|033|stroke-related inattention
C0233414|033|postictal inattention
C0233414|033|hypoxic attention deficit
C0233414|033|attention deficit – dementia
C0233414|033|vascular attention disturbance
C0233414|033|frontotemporal attention impairment
C0233414|033|alzheimer’s-related inattention
C0233414|033|pd-related inattention
C0233414|033|adhd (in context)
C0233414|033|cognitive slowing
C0233414|033|mental slowing
C0233414|033|bradyphrenia
C0233414|033|psychomotor slowing
C0233414|033|reduced cognitive speed
C0233414|033|attention lapses
C0233414|033|attentional lapses
C0233414|033|fluctuating loc with impaired attention
C0233414|033|impaired divided attention
C0233414|033|poor selective attention
C0233414|033|decreased sustained attention
C0233414|033|impaired sustained attention
C0233414|033|non-sustained attention
C0233414|033|poor task persistence
C0233414|033|vigilance deficit
C0233414|033|monitoring deficit
C0233414|033|reactivity impairment
C0233414|033|impaired responsiveness
C0233414|033|delayed responses
C0233414|033|slow to respond
C0233414|033|diminished alertness
C0233414|033|poor alertness
C0233414|033|reduced mental tracking
C0233414|033|errors in serial 7s
C0233414|033|errors on mmse attention
C0233414|033|failed world backward
C0233414|033|failed serial subtraction
C0233414|033|moca attention deficit
C0233414|033|mmse attention deficit
C0233414|033|consciousness disturbance
C0233414|033|consciousness fluctuation
C0233414|033|encephalopathic state
C0233414|033|encephalopathy with inattention
C0233414|033|cognitive disturbance
C0233414|033|attention-executive dysfunction
C0233414|033|difficulty following conversation
C0233414|033|easily dazed
C0233414|033|mentation fluctuating
C0233414|033|impaired cognitive control
C0233414|033|diffuse cognitive impairment
C0233414|033|loss of vigilance
C0233414|033|decreased mental flexibility
C0233414|033|reduced alertness and attention
C0233414|033|nonverbal inattention
C0233414|033|mild inattentiveness
C0233414|033|moderate inattentiveness
C0233414|033|severe inattentiveness
C0233414|033|attentional failures
C0233414|033|sustained concentration deficit
C0233414|033|task inattention
C0233414|033|slow processing speed
C0233414|033|difficulty maintaining attention
C0233414|033|difficulty with dual tasking
C0233414|033|attention span decreased
C0233414|033|slowed mentation
C0233414|033|impaired mental tracking
C0233414|033|errors on trail making
C0233414|033|omissions on attention tasks
C0233414|033|mental fatigue
C0233414|033|cognitive fatigue
C0233414|033|inattentive subtype
C0233414|033|inattentive presentation
C0454643|033|word finding difficulty
C0454643|033|word-finding difficulty
C0454643|033|word retrieval difficulty
C0454643|033|word finding disorder
C0454643|033|word-finding disorder
C0454643|033|word retrieval deficit
C0454643|033|word-finding deficit
C0454643|033|anomia
C0454643|033|anomic aphasia
C0454643|033|dysnomia
C0454643|033|dysnomia aphasia
C0454643|033|impaired word retrieval
C0454643|033|difficulty with naming
C0454643|033|naming deficit
C0454643|033|naming difficulty
C0454643|033|naming impairment
C0454643|033|impaired naming
C0454643|033|expressive anomia
C0454643|033|aphasia—anomic type
C0454643|033|aphasia (anomic)
C0454643|033|aphasic word-finding difficulty
C0454643|033|aphasic word finding
C0454643|033|aphasic dysnomia
C0454643|033|poststroke anomia
C0454643|033|ischemic anomia
C0454643|033|nonfluent anomia
C0454643|033|fluent anomia
C0454643|033|broca's aphasia with word-finding
C0454643|033|wernicke's aphasia with word-finding
C0454643|033|neurogenic anomia
C0454643|033|vascular anomia
C0454643|033|dementia-related anomia
C0454643|033|ad anomia
C0454643|033|alzheimer's related anomia
C0454643|033|ftd anomia
C0454643|033|semantic anomia
C0454643|033|progressive anomia
C0454643|033|ppa anomia
C0454643|033|primary progressive aphasia with anomia
C0454643|033|tbi-related word-finding
C0454643|033|chemo-induced anomia
C0454643|033|postictal word-finding
C0454643|033|migraine-related word-finding
C0454643|033|tia-related word-finding
C0454643|033|transient anomia
C0454643|033|acute anomia
C0454643|033|chronic anomia
C0454643|033|receptive anomia
C0454643|033|expressive dysnomia
C0454643|033|mild anomic aphasia
C0454643|033|mild word-finding deficit
C0454643|033|moderate word-finding deficit
C0454643|033|severe word-finding impairment
C0454643|033|anomic type aphasia
C0454643|033|amnestic aphasia
C0454643|033|loc anomia
C0454643|033|post-op word-finding
C0454643|033|perseverative anomia
C0454643|033|lexical retrieval deficit
C0454643|033|word retrieval impairment
C0454643|033|verbal retrieval deficit
C0454643|033|verbal retrieval impairment
C0454643|033|verbal anomia
C0454643|033|language retrieval deficit
C0454643|033|language retrieval difficulty
C0454643|033|tip-of-the-tongue state
C0454643|033|tot phenomenon
C0454643|033|speech output deficit
C0454643|033|speech hesitation
C0454643|033|lexical-access deficit
C0454643|033|semantic retrieval deficit
C0454643|033|lexical access disorder
C0454643|033|naming latency
C0454643|033|naming hesitation
C0454643|033|naming block
C0454643|033|repetitive anomic errors
C0454643|033|searching for words
C0454643|033|circumlocutory speech
C0454643|033|circumlocution due to anomia
C0454643|033|paraphasic naming errors
C0454643|033|semantic paraphasia (word-finding)
C0454643|033|phonemic paraphasia (word-finding)
C0454643|033|word-finding pauses
C0454643|033|speech arrest (anomia)
C0454643|033|motor aphasia—anomic
C0454643|033|nonfluent aphasia with anomia
C0454643|033|fluent aphasia with anomia
C0454643|033|thalamic anomia
C0454643|033|broca-type word-finding
C0454643|033|wernicke-type word-finding
C0454643|033|global aphasia (with word-finding)
C0454643|033|pca-related anomia
C0454643|033|temporal lobe anomia
C0454643|033|parietal lobe anomia
C0454643|033|frontal lobe anomia
C0454643|033|multifactorial anomia
C0454643|033|amnestic speech
C0454643|033|amnestic disorder with aphasia
C0454643|033|unclassifiable aphasia—anomia dominant
C0454643|033|lbd-related anomia
C0454643|033|vad anomia
C0454643|033|cva anomia
C0454643|033|stroke-related anomia
C0454643|033|sah-related anomia
C0454643|033|functional word-finding
C0454643|033|functional anomia
C0454643|033|psychogenic word-finding issues
C0454643|033|depression-related anomia
C0454643|033|delirium-associated anomia
C0454643|033|delirium word-finding
C0454643|033|focal word-finding deficit
C0454643|033|transient expressive aphasia
C0454643|033|transient expressive anomia
C0454643|033|mild cognitive impairment with anomia
C0454643|033|mci anomia
C0454643|033|age-related word-finding
C0454643|033|developmental anomia
C0454643|033|childhood anomia
C0454643|033|congenital anomia
C0454643|033|genetic anomia
C0454643|033|drug-induced anomia
C0454643|033|medication-induced anomia
C0454643|033|toxic-metabolic word-finding
C0454643|033|metabolic anomia
C0454643|033|encephalopathic anomia
C0454643|033|encephalopathy word-finding
C0454643|033|post-concussive word-finding
C0454643|033|remote word-finding deficit
C0454643|033|hypertensive word-finding
C0454643|033|amyloid anomia
C0454643|033|infectious aphasia—anomic
C0454643|033|autoimmune anomia
C0454643|033|paraneoplastic anomia
C0454643|033|radiation-induced anomia
C0454643|033|postradiation word-finding
C0454643|033|paraphasic speech (anomia)
C0454643|033|mixed aphasia with anomia
C0454643|033|multilingual anomia
C0454643|033|multilingual naming deficit
C0454643|033|secondary anomia
C0454643|033|primary anomia
C0454643|033|acquired anomia
C0454643|033|post-traumatic anomia
C0454643|033|postinfectious word-finding
C0454643|033|postencephalitic anomia
C0454643|033|retograde anomia
C0454643|033|anomic variant ppa
C0454643|033|semantic variant ppa
C0454643|033|logopenic variant ppa with anomia
C0454643|033|logopenic word-finding
C0454643|033|speech disruption (anomic)
C0454643|033|speech disturbance—anomia
C0454643|033|language disturbance—anomia
C0454643|033|pragmatic anomia
C0454643|033|compensated anomia
C0454643|033|residual aphasia—anomic
C0454643|033|remitted aphasia—anomic
C0454643|033|active word-finding deficit
C0454643|033|intermittent word-finding
C0454643|033|cathartic anomia
C0454643|033|verbal access disorder
C0454643|033|lexical semantic deficit
C0454643|033|impaired expressive language (naming)
C0454643|033|aphasia nos (anomic features)
C0454643|033|word-finding issue
C0454643|033|naming problem
C0542476|033|forgetful
C0542476|033|forgetfulness
C0542476|033|memory loss
C0542476|033|memory impairment
C0542476|033|impaired memory
C0542476|033|amnesia
C0542476|033|amnesic
C0542476|033|dementia
C0542476|033|cognitive decline
C0542476|033|cognitive impairment
C0542476|033|dec cognition
C0542476|033|dec memory
C0542476|033|declining memory
C0542476|033|short-term memory loss
C0542476|033|impaired recall
C0542476|033|poor recall
C0542476|033|dec recall
C0542476|033|difficulty remembering
C0542476|033|difficulty recalling
C0542476|033|absent-minded
C0542476|033|absentmindedness
C0542476|033|lapses in memory
C0542476|033|slips of memory
C0542476|033|confused
C0542476|033|confusion
C0542476|033|mental fog
C0542476|033|mentally foggy
C0542476|033|disoriented
C0542476|033|disorientation
C0542476|033|impaired recent memory
C0542476|033|imp rec mem
C0542476|033|impaired remote memory
C0542476|033|imp rem mem
C0542476|033|anterograde amnesia
C0542476|033|retrograde amnesia
C0542476|033|transient global amnesia
C0542476|033|mnestic deficit
C0542476|033|mnemonic deficit
C0542476|033|forgetting
C0542476|033|trouble remembering
C0542476|033|trouble recalling
C0542476|033|trouble with memory
C0542476|033|stms loss
C0542476|033|ltms loss
C0542476|033|short-term mem loss
C0542476|033|long-term mem loss
C0542476|033|impaired working memory
C0542476|033|deficits in memory
C0542476|033|executive dysfunction
C0542476|033|mild cognitive impairment
C0542476|033|mci
C0542476|033|early dementia
C0542476|033|alzheimer's type memory loss
C0542476|033|ad-type memory loss
C0542476|033|vascular memory impairment
C0542476|033|vascular cognitive impairment
C0542476|033|post-stroke memory loss
C0542476|033|stroke-related memory loss
C0542476|033|ischemic memory loss
C0542476|033|tbi-related memory loss
C0542476|033|trauma-induced amnesia
C0542476|033|chemobrain
C0542476|033|chemo-induced cognitive impairment
C0542476|033|chemo-induced memory loss
C0542476|033|delirium
C0542476|033|encephalopathic
C0542476|033|encephalopathy-related memory loss
C0542476|033|hiv-associated neurocognitive disorder
C0542476|033|metabolic memory impairment
C0542476|033|hepatic encephalopathy memory loss
C0542476|033|alcohol-related memory loss
C0542476|033|korsakoff syndrome
C0542476|033|wernicke-korsakoff
C0542476|033|anoxic memory loss
C0542476|033|hypoxic memory loss
C0542476|033|hypoglycemia-related memory loss
C0542476|033|thyroid-related memory impairment
C0542476|033|hypothyroid memory loss
C0542476|033|aging-related memory loss
C0542476|033|age-assoc memory change
C0542476|033|age-assoc mem loss
C0542476|033|senile memory impairment
C0542476|033|senile forgetfulness
C0542476|033|senile dementia
C0542476|033|lewy body-related memory loss
C0542476|033|dlb-associated memory impairment
C0542476|033|frontotemporal memory loss
C0542476|033|ftd-associated memory impairment
C0542476|033|parkinsonian memory impairment
C0542476|033|parkinson's-related memory loss
C0542476|033|pd-associated memory impairment
C0542476|033|ms-related memory impairment
C0542476|033|multiple sclerosis memory loss
C0542476|033|amnestic
C0542476|033|cbi (cognitive behavioral impairment)
C0542476|033|intellectual decline
C0542476|033|progressive memory loss
C0542476|033|transient memory loss
C0542476|033|forgetting names
C0542476|033|forgetting appointments
C0542476|033|repeat questioning
C0542476|033|losing items
C0542476|033|difficulty learning new info
C0542476|033|dysmnestic
C0542476|033|declining cognition
C0542476|033|impaired recognition
C0542476|033|impaired information retention
C0542476|033|impaired learning
C0542476|033|forgetfulness episodes
C0542476|033|episodic memory loss
C0542476|033|impaired autobiographical memory
C0542476|033|poor memory
C0542476|033|dec memory retention
C0542476|033|deficient memory
C0542476|033|suboptimal memory
C0542476|033|slowed mental processing
C0542476|033|impairment in recall
C0542476|033|impaired recent recall
C0542476|033|impaired delayed recall
C0542476|033|inconsistent recall
C0542476|033|diminished memory capacity
C0542476|033|lapses in recall
C0542476|033|poor retention
C0542476|033|memory difficulties
C0542476|033|problems with memory
C0542476|033|diminished short-term memory
C0542476|033|lack of recall
C0542476|033|absent recall
C0542476|033|frontal lobe memory impairment
C0542476|033|temporal lobe memory impairment
C0542476|033|difficulty storing new memories
C0542476|033|working memory difficulty
C0542476|033|amnesia nos
C0542476|033|cognitive deficits
C0542476|033|short term memory impairment
C0542476|033|long term memory impairment
C0542476|033|decline in stm
C0542476|033|decline in ltm
C0542476|033|stm impairment
C0542476|033|ltm impairment
C0542476|033|frequent forgetting
C0542476|033|recurrent memory lapses
C0542476|033|frequent memory lapses
C0542476|033|decreased new learning
C0542476|033|impaired ability to recall facts
C0542476|033|hippocampal memory loss
C0542476|033|executive memory dysfunction
C0542476|033|amnesic episode
C0542476|033|mnestic disturbance
C0542476|033|forgets instructions
C0542476|033|forgetting conversations
C0542476|033|disrupted memory
C0542476|033|amnesic disorder
C0542476|033|amnesic syndrome
C0542476|033|impaired consolidation
C0542476|033|delayed retrieval
C0542476|033|impaired encoding
C0542476|033|imp encoding
C0542476|033|imp retrieval
C0542476|033|impaired retrieval
C1522449|061|radiation therapy
C1522449|061|radiotherapy
C1522449|061|rt
C1522449|061|xrt
C1522449|061|external beam radiation
C1522449|061|external beam rt
C1522449|061|external beam radiotherapy
C1522449|061|ebrt
C1522449|061|radiation tx
C1522449|061|rad tx
C1522449|061|rad therapy
C1522449|061|radio tx
C1522449|061|ionizing radiation therapy
C1522449|061|therapeutic irradiation
C1522449|061|irradiation
C1522449|061|radiotherapeutic procedure
C1522449|061|radiotherapeutics
C1522449|061|radioisotope therapy
C1522449|061|teletherapy
C1522449|061|brachytherapy
C1522449|061|imrt
C1522449|061|intensity-modulated rt
C1522449|061|intensity-modulated radiation therapy
C1522449|061|igrt
C1522449|061|image-guided radiation therapy
C1522449|061|stereotactic radiosurgery
C1522449|061|srs
C1522449|061|sbrt
C1522449|061|stereotactic body radiation therapy
C1522449|061|proton therapy
C1522449|061|proton beam therapy
C1522449|061|pbt
C1522449|061|conventional radiation
C1522449|061|fractionated radiation
C1522449|061|adjuvant rt
C1522449|061|neoadjuvant rt
C1522449|061|conformal rt
C1522449|061|3d crt
C1522449|061|3d conformal radiation
C1522449|061|3d conformal rt
C1522449|061|three-dimensional conformal rt
C1522449|061|pall rt
C1522449|061|palliative radiation
C1522449|061|palliative rt
C1522449|061|whole brain rt
C1522449|061|cns rt
C1522449|061|cranial radiation
C1522449|061|tbi
C1522449|061|total body irradiation
C1522449|061|prophylactic cranial irradiation
C1522449|061|pci
C1522449|061|accelerated rt
C1522449|061|boost radiation
C1522449|061|boost rt
C1522449|061|intraoperative rt
C1522449|061|iort
C1522449|061|rad onc tx
C1522449|061|rad oncology therapy
C1522449|061|radiation course
C1522449|061|external radiation
C1522449|061|radiation
C1522450|061|brachy
C1522451|061|intraop rt
C1522452|061|intraop radiation
C1522453|061|wbrt
C1522454|061|srt
C1522455|061|radiosurgery
C1522456|061|proton
C1522457|061|electron
C1522458|061|photon
C1522459|061|vmat
C1522460|061|volumetric modulated arc radiotherapy
