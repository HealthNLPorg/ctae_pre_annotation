C0018801|000|heart failure
C0018801|000|hf
C0018801|000|congestive heart failure
C0018801|000|chf
C0018801|000|acute heart failure
C0018801|000|acute hf
C0018801|000|chronic heart failure
C0018801|000|chronic hf
C0018801|000|decompensated heart failure
C0018801|000|decompensated hf
C0018801|000|compensated heart failure
C0018801|000|compensated hf
C0018801|000|high-output heart failure
C0018801|000|hof
C0018801|000|low-output heart failure
C0018801|000|lof
C0018801|000|right heart failure
C0018801|000|right-sided heart failure
C0018801|000|right hf
C0018801|000|left heart failure
C0018801|000|left-sided heart failure
C0018801|000|left hf
C0018801|000|biventricular heart failure
C0018801|000|biventricular hf
C0018801|000|diastolic heart failure
C0018801|000|dhf
C0018801|000|heart failure with preserved ejection fraction
C0018801|000|hfpef
C0018801|000|preserved ef heart failure
C0018801|000|systolic heart failure
C0018801|000|shf
C0018801|000|heart failure with reduced ejection fraction
C0018801|000|hfref
C0018801|000|reduced ef heart failure
C0018801|000|borderline ef heart failure
C0018801|000|mid-range ef heart failure
C0018801|000|hfmref
C0018801|000|ischemic heart failure
C0018801|000|ischemic hf
C0018801|000|nonischemic heart failure
C0018801|000|nonischemic hf
C0018801|000|valvular heart failure
C0018801|000|valvular hf
C0018801|000|hypertensive heart failure
C0018801|000|hypertensive hf
C0018801|000|amyloid heart failure
C0018801|000|amyloidosis-related hf
C0018801|000|cardiac amyloidosis with failure
C0018801|000|chemotherapy-induced heart failure
C0018801|000|chemo-induced hf
C0018801|000|ppcm
C0018801|000|peripartum cardiomyopathy
C0018801|000|tachycardia-induced heart failure
C0018801|000|tachycardia-induced hf
C0018801|000|myocarditis-induced heart failure
C0018801|000|myocarditis-related hf
C0018801|000|alcoholic cardiomyopathy with failure
C0018801|000|alcohol-related heart failure
C0018801|000|infiltrative cardiomyopathy with failure
C0018801|000|viral cardiomyopathy with failure
C0018801|000|postpartum heart failure
C0018801|000|dilated cardiomyopathy with failure
C0018801|000|dilated cm with hf
C0018801|000|idiopathic heart failure
C0018801|000|familial heart failure
C0018801|000|restrictive cardiomyopathy with failure
C0018801|000|rcm with hf
C0018801|000|cardiomyopathy with failure
C0018801|000|cm with hf
C0018801|000|advanced heart failure
C0018801|000|end-stage heart failure
C0018801|000|terminal heart failure
C0018801|000|refractory heart failure
C0018801|000|progressive heart failure
C0018801|000|acute on chronic heart failure
C0018801|000|aoc heart failure
C0018801|000|post-mi heart failure
C0018801|000|post-infarction heart failure
C0018801|000|cardiorenal syndrome
C0018801|000|crs
C0018801|000|pulmonary edema due to chf
C0018801|000|pump failure
C0018801|000|cardiac failure
C0018801|000|ventricular failure
C0018801|000|ventricular dysfunction
C0018801|000|lv failure
C0018801|000|left ventricular failure
C0018801|000|rv failure
C0018801|000|right ventricular failure
C0018801|000|congestive cardiac failure
C0018801|000|ccf
C0018801|000|preload failure
C0018801|000|forward failure
C0018801|000|backward failure
C0018801|000|cardiac decompensation
C0018801|000|volume overload chf
C0018801|000|volume overload hf
C0018801|000|fluid overload chf
C0018801|000|fluid overload hf
C0018801|000|exacerbated chf
C0018801|000|exacerbation of hf
C0018801|000|cardiogenic pulmonary edema
C0018801|000|pulmonary congestion due to hf
C0018801|000|post-cardiac surgery hf
C0018801|000|iatrogenic heart failure
C0018801|000|drug-induced heart failure
C0018801|000|radiation-induced heart failure
C0018801|000|cor pulmonale with failure
C0018801|000|cor pulmonale with chf
C0018801|000|secondary heart failure
C0018801|000|primary heart failure
C0018801|000|tachyarrhythmia-related heart failure
C0018801|000|bradycardia-induced heart failure
C0018801|000|hfref exacerbation
C0018801|000|hfpef exacerbation
C0018801|000|heart failure with mid-range ef
C0018801|000|heart failure with mildly reduced ef
C0018801|000|diabetic cardiomyopathy with failure
C0018801|000|dm-related heart failure
C0018801|000|obesity-related heart failure
C0018801|000|thyrotoxic heart failure
C0018801|000|thyroid disease–related hf
C0018801|000|constrictive pericarditis with failure
C0018801|000|volume overloaded heart
C0018801|000|chf exacerbation
C0018801|000|new-onset heart failure
C0018801|000|new hf
C0018801|000|acute decompensated heart failure
C0018801|000|adhf
C0018801|000|cardiac insufficiency
C0018801|000|chronic decompensated heart failure
C0018801|000|acute exacerbation of chf
C0018801|000|exertional heart failure
C0018801|000|post-viral heart failure
C0018801|000|post-viral cardiomyopathy with failure
C0018801|000|pericardial disease with failure
C0018801|000|transfusion-associated circulatory overload
C0018801|000|taco
C0018801|000|heart failure secondary to anemia
C0018801|000|high-output cardiac failure
C0018801|000|myocardial failure
C0018801|000|congestive myocardial failure
C0018801|000|acute left ventricular failure
C0018801|000|acute lvf
C0018801|000|chronic right heart failure
C0018801|000|heart failure with arrhythmia
C0018801|000|arrhythmia-related heart failure
C0018801|000|post-cardiotomy heart failure
C0018801|000|post-transplant heart failure
C0018801|000|transplant heart failure
C0018801|000|device-related heart failure
C0018801|000|lvad-related hf
C0018801|000|right heart dysfunction
C0018801|000|left heart dysfunction
C0018801|000|cardiac pump failure
C0018801|000|post-ischemic heart failure
C0018801|000|ischemic dilated cardiomyopathy with failure
C0018801|000|post-reperfusion heart failure
C0018801|000|stress-induced cardiomyopathy with failure
C0018801|000|takotsubo with failure
C0018801|000|takotsubo hf
C0018801|000|chagas disease with heart failure
C0018801|000|hereditary heart failure
C0018801|000|arvc with failure
C0018801|000|arrhythmogenic rv cardiomyopathy with hf
C0027051|000|myocardial infarction
C0027051|000|mi
C0027051|000|acute mi
C0027051|000|ami
C0027051|000|acute myocardial infarction
C0027051|000|stemi
C0027051|000|st-elevation mi
C0027051|000|st-elevation myocardial infarction
C0027051|000|nstemi
C0027051|000|non-st-elevation mi
C0027051|000|non-st-elevation myocardial infarction
C0027051|000|transmural mi
C0027051|000|subendocardial mi
C0027051|000|inferior mi
C0027051|000|anterior mi
C0027051|000|lateral mi
C0027051|000|posterior mi
C0027051|000|septal mi
C0027051|000|high lateral mi
C0027051|000|unstable coronary syndrome
C0027051|000|ischemic mi
C0027051|000|ischemic infarct
C0027051|000|cardiac infarct
C0027051|000|acute coronary syndrome
C0027051|000|acs
C0027051|000|coronary thrombosis
C0027051|000|coronary occlusion
C0027051|000|transmural infarct
C0027051|000|subendocardial infarct
C0027051|000|heart attack
C0027051|000|old mi
C0027051|000|prior mi
C0027051|000|healed mi
C0027051|000|silent infarction
C0027051|000|silent mi
C0027051|000|q wave mi
C0027051|000|non-q wave mi
C0027051|000|spontaneous mi
C0027051|000|type 1 mi
C0027051|000|type i mi
C0027051|000|type 2 mi
C0027051|000|type ii mi
C0027051|000|demand mi
C0027051|000|supply-demand mismatch mi
C0027051|000|secondary mi
C0027051|000|perioperative mi
C0027051|000|post-procedure mi
C0027051|000|stent thrombosis mi
C0027051|000|in-stent mi
C0027051|000|valvular mi
C0027051|000|hypertensive mi
C0027051|000|amyloid mi
C0027051|000|chemo-induced mi
C0027051|000|cancer therapy–related mi
C0027051|000|ppcm-related mi
C0027051|000|post-partum cm with mi
C0027051|000|myocarditis-related mi
C0027051|000|tachycardia-induced mi
C0027051|000|atrial fibrillation mi
C0027051|000|coronary embolism mi
C0027051|000|embolism-related mi
C0027051|000|coronary spasm mi
C0027051|000|vasospastic mi
C0027051|000|coronary dissection mi
C0027051|000|scad mi
C0027051|000|spontaneous coronary artery dissection mi
C0027051|000|thrombotic mi
C0027051|000|microvascular mi
C0027051|000|microvascular infarction
C0027051|000|cardiac necrosis
C0027051|000|myocardial necrosis
C0027051|000|myocardial injury (ischemic)
C0027051|000|ischemia-induced necrosis
C0027051|000|supply-demand mismatch infarct
C0027051|000|lv infarct
C0027051|000|rv infarct
C0027051|000|presumed mi
C0027051|000|possible mi
C0027051|000|probable mi
C0027051|000|unrecognized mi
C0027051|000|nontransmural mi
C0027051|000|recurrent mi
C0027051|000|multiple mi
C0027051|000|re-infarction
C0027051|000|reinfarction
C0027051|000|reinfarct
C0027051|000|reinfarcted myocardium
C0027051|000|extensive mi
C0027051|000|widespread mi
C0027051|000|limited mi
C0027051|000|microscopic mi
C0027051|000|multi-territory mi
C0027051|000|multivessel mi
C0027051|000|single vessel mi
C0027051|000|inferolateral mi
C0027051|000|anterolateral mi
C0027051|000|posterolateral mi
C0027051|000|apical mi
C0027051|000|basal mi
C0027051|000|old inferior mi
C0027051|000|old anterior mi
C0027051|000|old lateral mi
C0027051|000|old septal mi
C0027051|000|old transmural mi
C0027051|000|old subendocardial mi
C0027051|000|silent anterior mi
C0027051|000|silent inferior mi
C0027051|000|silent posterior mi
C0027051|000|acute infarct
C0027051|000|acute transmural mi
C0027051|000|acute subendocardial mi
C0027051|000|acute anterior mi
C0027051|000|acute inferior mi
C0027051|000|acute lateral mi
C0027051|000|acute septal mi
C0027051|000|acute posterior mi
C0027051|000|nstemi acs
C0027051|000|stemi acs
C0027051|000|post-cath mi
C0027051|000|periprocedural mi
C0027051|000|high sensitivity troponin mi
C0027051|000|troponin-positive mi
C0027051|000|troponin rise (mi)
C0027051|000|ihd with mi
C0027051|000|ischemic heart disease with mi
C0027051|000|cad with mi
C0027051|000|coronary artery disease with mi
C0027051|000|mi with lv dysfunction
C0027051|000|mi with heart failure
C0027051|000|chf secondary to mi
C0027051|000|ventricular infarct
C0027051|000|coronary syndrome (mi)
C0027051|000|infarcted myocardium
C0027051|000|myocardial infarct tissue
C0027051|000|fibrotic myocardium post mi
C0027051|000|scarred myocardium (post mi)
C0027051|000|cardiac event (infarct)
C0027051|000|myocardial event (inf. type)
C0027051|000|myocardial ischemia with infarction
C0027051|000|ischemic cardiomyopathy (mi)
C0027051|000|mi secondary to embolus
C0027051|000|mi secondary to spasm
C0027051|000|mi secondary to amyloid
C0027051|000|mi secondary to hypotension
C0027051|000|mi secondary to vasospasm
C0027051|000|mi secondary to thrombosis
C0027051|000|mi secondary to hypertension
C0027051|000|mi secondary to cocaine
C0027051|000|cocaine-induced mi
C0027051|000|mi secondary to anemia
C0027051|000|demand ischemia with infarct
C0027051|000|coronary supply mi
C0027051|000|coronary demand mi
C0027051|000|type 3 mi
C0027051|000|type iii mi
C0027051|000|type 4a mi
C0027051|000|type 4b mi
C0027051|000|type 4c mi
C0027051|000|type 5 mi
C0027051|000|post-pci mi
C0027051|000|post-cabg mi
C0027051|000|late mi
C0027051|000|early mi
C0027051|000|periinfarct
C0027051|000|myocardial infarct zone
C0027051|000|mi territory
C0027051|000|coronary syndrome (with mi)
C0027051|000|infarct-related artery
C0027051|000|culprit lesion mi
C0027051|000|mi with papillary muscle involvement
C0027051|000|acute infarction event
C0027051|000|cardiac event (mi type)
C0027051|000|coronary syndrome with infarct
C0027051|000|cardiac ischemic event
C0027051|000|acute plaque rupture mi
C0027051|000|mi with thrombus
C0002965|000|unstable angina
C0002965|000|ua
C0002965|000|usa
C0002965|000|acs-ua
C0002965|000|pre-infarction angina
C0002965|000|crescendo angina
C0002965|000|intermediate coronary syndrome
C0002965|000|preinfarction angina
C0002965|000|threatened mi
C0002965|000|angina at rest
C0002965|000|rest angina
C0002965|000|ischemic ua
C0002965|000|ischemic unstable angina
C0002965|000|acute isch angina
C0002965|000|non-st elevation acs-ua
C0002965|000|nstemi/ua
C0002965|000|nstemi rule out
C0002965|000|nstemi suspected/ua
C0002965|000|decubitus ua
C0002965|000|variant ua
C0002965|000|refractory ua
C0002965|000|angina exacerbation
C0002965|000|progressive angina
C0002965|000|worsening angina
C0002965|000|dynamic angina
C0002965|000|unstable exertional angina
C0002965|000|secondary unstable angina
C0002965|000|valvular ua
C0002965|000|valvular unstable angina
C0002965|000|hypertensive ua
C0002965|000|hypertensive unstable angina
C0002965|000|chemo-induced unstable angina
C0002965|000|drug-induced ua
C0002965|000|myocarditis-associated ua
C0002965|000|tachycardia-induced ua
C0002965|000|ppcm with ua
C0002965|000|nonischemic ua
C0002965|000|postintervention ua
C0002965|000|post-pci ua
C0002965|000|post-cabg ua
C0002965|000|bypass ua
C0002965|000|stent ua
C0002965|000|spontaneous unstable angina
C0002965|000|recurrent ua
C0002965|000|recurring unstable angina
C0002965|000|intractable ua
C0002965|000|resistant unstable angina
C0002965|000|unstable post-infarct angina
C0002965|000|angina instable
C0002965|000|instable angina
C0002965|000|angor instable
C0002965|000|ua/nstemi
C0002965|000|non-q-wave ua
C0002965|000|noq ua
C0002965|000|unstable ep angina
C0002965|000|ua w/elevated troponin
C0002965|000|ua (tn-)
C0038454|000|cerebrovascular accident
C0038454|000|cva
C0038454|000|stroke
C0038454|000|acute stroke
C0038454|000|embolic stroke
C0038454|000|thrombotic stroke
C0038454|000|hemorrhagic stroke
C0038454|000|ischemic stroke
C0038454|000|nonischemic stroke
C0038454|000|lacunar stroke
C0038454|000|cerebral infarct
C0038454|000|cerebral infarction
C0038454|000|cerebral hemorrhage
C0038454|000|brain attack
C0038454|000|brain infarct
C0038454|000|brain infarction
C0038454|000|acute cerebral infarct
C0038454|000|large vessel stroke
C0038454|000|small vessel stroke
C0038454|000|cryptogenic stroke
C0038454|000|watershed infarct
C0038454|000|tia with infarct
C0038454|000|intraparenchymal hemorrhage
C0038454|000|parenchymal hemorrhage
C0038454|000|icvh
C0038454|000|ich
C0038454|000|intracerebral hemorrhage
C0038454|000|subcortical infarct
C0038454|000|cortical infarct
C0038454|000|pca stroke
C0038454|000|mca stroke
C0038454|000|aca stroke
C0038454|000|posterior stroke
C0038454|000|anterior circulation stroke
C0038454|000|posterior circulation stroke
C0038454|000|valvular embolic stroke
C0038454|000|cardioembolic stroke
C0038454|000|atrial fib stroke
C0038454|000|afib stroke
C0038454|000|non-valvular stroke
C0038454|000|artery-to-artery embolic stroke
C0038454|000|arterial embolic stroke
C0038454|000|vertebrobasilar stroke
C0038454|000|basilar stroke
C0038454|000|brainstem stroke
C0038454|000|pontine stroke
C0038454|000|cerebellar stroke
C0038454|000|subarachnoid hemorrhage
C0038454|000|sah
C0038454|000|midline cerebral infarct
C0038454|000|right mca stroke
C0038454|000|left mca stroke
C0038454|000|r mca infarct
C0038454|000|l mca infarct
C0038454|000|left hemisphere infarct
C0038454|000|right hemisphere infarct
C0038454|000|r cortical stroke
C0038454|000|l cortical stroke
C0038454|000|chronic infarct
C0038454|000|acute on chronic infarct
C0038454|000|microvascular infarct
C0038454|000|silent infarct
C0038454|000|old infarct
C0038454|000|remote infarct
C0038454|000|multi-infarct
C0038454|000|multiple infarcts
C0038454|000|multi-territorial stroke
C0038454|000|transient cerebral ischemia
C0038454|000|cerebral ischemia
C0038454|000|acute cerebral ischemia
C0038454|000|territorial infarct
C0038454|000|territorial stroke
C0038454|000|territorial hemorrhage
C0038454|000|flow-related infarct
C0038454|000|global cerebral ischemia
C0038454|000|atherothrombotic stroke
C0038454|000|cholesterol embolic stroke
C0038454|000|calcific embolic stroke
C0038454|000|infective embolic stroke
C0038454|000|meningovascular stroke
C0038454|000|arteriopathic stroke
C0038454|000|hypertensive stroke
C0038454|000|hypertensive intracerebral hemorrhage
C0038454|000|amyloid angiopathy stroke
C0038454|000|amyloid angiopathy hemorrhage
C0038454|000|caa-associated hemorrhage
C0038454|000|leukoaraiosis-associated stroke
C0038454|000|chemo-induced stroke
C0038454|000|radiation-induced stroke
C0038454|000|drug-induced stroke
C0038454|000|ppcm-related stroke
C0038454|000|peripartum stroke
C0038454|000|pregnancy-associated stroke
C0038454|000|puerperal stroke
C0038454|000|myocarditis-associated stroke
C0038454|000|tachycardia-induced stroke
C0038454|000|arrhythmic embolic stroke
C0038454|000|endocarditis embolic stroke
C0038454|000|paradoxical embolic stroke
C0038454|000|nonbacterial thrombotic embolic stroke
C0038454|000|nbte stroke
C0038454|000|moya moya stroke
C0038454|000|vasculitis-associated stroke
C0038454|000|sle-associated stroke
C0038454|000|antiphospholipid stroke
C0038454|000|hypercoagulable stroke
C0038454|000|coagulopathy stroke
C0038454|000|cocaine-induced stroke
C0038454|000|vasospasm-associated infarct
C0038454|000|hypoperfusion stroke
C0038454|000|hemodynamic stroke
C0038454|000|low-flow infarct
C0038454|000|occlusive stroke
C0038454|000|arterial occlusive infarct
C0038454|000|arterial occlusion stroke
C0038454|000|large artery atherosclerotic stroke
C0038454|000|laa stroke
C0038454|000|intracranial atherosclerotic stroke
C0038454|000|extracranial atherosclerotic stroke
C0038454|000|atherothrombotic infarct
C0038454|000|cavitary infarct
C0038454|000|cavitating infarct
C0038454|000|encephalomalacic infarct
C0038454|000|encephalomalacia from cva
C0038454|000|cerebellar infarct
C0038454|000|cerebellar hemorrhage
C0038454|000|medullary infarct
C0038454|000|medullary stroke
C0038454|000|brainstem infarct
C0038454|000|thalamic infarct
C0038454|000|thalamic hemorrhage
C0038454|000|putaminal hemorrhage
C0038454|000|putaminal infarct
C0038454|000|capsular stroke
C0038454|000|internal capsule infarct
C0038454|000|subcortical hemorrhage
C0038454|000|subcortical stroke
C0038454|000|watershed stroke
C0038454|000|borderzone infarct
C0038454|000|lacunar infarct
C0038454|000|peri-ictal infarct
C0038454|000|hypoxic ischemic stroke
C0038454|000|cardiac arrest-related stroke
C0038454|000|post-cardiac arrest infarct
C0038454|000|cerebral embolism
C0038454|000|cerebral embolic event
C0038454|000|cerebral thromboembolism
C0038454|000|cerebrovascular event
C0038454|000|acute cerebrovascular event
C0038454|000|major stroke
C0038454|000|minor stroke
C0038454|000|silent stroke
C0038454|000|subclinical stroke
C0038454|000|cerebral event
C0038454|000|pres-associated infarct
C0038454|000|posterior reversible encephalopathy stroke
C0038454|000|arteriopathy-associated infarct
C0038454|000|cortical laminar necrosis
C0038454|000|subdural hematoma stroke
C0038454|000|cortical microinfarct
C0038454|000|cortical microbleed associated stroke
C0038454|000|embolism to brain
C0038454|000|embolus to brain
C0038454|000|cerebral occlusion event
C0038454|000|cerebral arterial infarct
C0038454|000|cerebral embologenic event
C0038454|000|left hemispheric stroke
C0038454|000|right hemispheric stroke
C0038454|000|left parietal stroke
C0038454|000|right parietal stroke
C0038454|000|left frontal infarct
C0038454|000|right frontal infarct
C0004238|000|atrial fibrillation
C0004238|000|af
C0004238|000|afib
C0004238|000|a-fib
C0004238|000|a fibrillation
C0004238|000|chronic atrial fibrillation
C0004238|000|paroxysmal atrial fibrillation
C0004238|000|persistent atrial fibrillation
C0004238|000|permanent atrial fibrillation
C0004238|000|long-standing persistent atrial fibrillation
C0004238|000|valvular atrial fibrillation
C0004238|000|nonvalvular atrial fibrillation
C0004238|000|nvaf
C0004238|000|valvular af
C0004238|000|nonvalvular af
C0004238|000|secondary atrial fibrillation
C0004238|000|recurrent atrial fibrillation
C0004238|000|acute atrial fibrillation
C0004238|000|postoperative atrial fibrillation
C0004238|000|poaf
C0004238|000|new-onset atrial fibrillation
C0004238|000|lone atrial fibrillation
C0004238|000|ischemic atrial fibrillation
C0004238|000|nonischemic atrial fibrillation
C0004238|000|hypertensive atrial fibrillation
C0004238|000|amyloid atrial fibrillation
C0004238|000|amyloidosis-related af
C0004238|000|chemo-induced atrial fibrillation
C0004238|000|chemotherapy-related af
C0004238|000|tachycardia-induced atrial fibrillation
C0004238|000|tachy-induced af
C0004238|000|ppcm-related atrial fibrillation
C0004238|000|peripartum af
C0004238|000|myocarditis-associated af
C0004238|000|alcoholic af
C0004238|000|holiday heart syndrome
C0004238|000|alcohol-induced atrial fibrillation
C0004238|000|af with rvr
C0004238|000|atrial fibrillation with rapid ventricular response
C0004238|000|af w/ rvr
C0004238|000|af with slow ventricular response
C0004238|000|af with bradycardia
C0004238|000|subclinical atrial fibrillation
C0004238|000|asymptomatic atrial fibrillation
C0004238|000|symptomatic atrial fibrillation
C0004238|000|atrial fib
C0004238|000|atrial-fib
C0004238|000|fib/flutter
C0004238|000|af/flutter
C0004238|000|af/afl
C0004238|000|a fib/flutter
C0004238|000|paroxysmal af
C0004238|000|persistent af
C0004238|000|permanent af
C0004238|000|long-standing persistent af
C0004238|000|recurrent af
C0004238|000|secondary af
C0004238|000|acute af
C0004238|000|new-onset af
C0004238|000|postop af
C0004238|000|post-op af
C0004238|000|common-type atrial fibrillation
C0004238|000|rapid atrial fibrillation
C0004238|000|atrial fibrillation crisis
C0004238|000|resistant atrial fibrillation
C0004238|000|uncontrolled atrial fibrillation
C0004238|000|controlled atrial fibrillation
C0004238|000|atf
C0004238|000|a. fib.
C0004238|000|a/f
C0004238|000|a-fibrillation
C0004238|000|afib p/w rvr
C0004238|000|paroxysmal a-fib
C0004238|000|persistent a-fib
C0004238|000|permanent a-fib
C0004238|000|af with slow vr
C0004238|000|af w/ svr
C0004238|000|valvular a-fib
C0004238|000|nonvalvular a-fib
C0004238|000|non-ischemic af
C0004238|000|ischemic af
C0004238|000|hypertensive af
C0004238|000|ms/af
C0004238|000|mitral stenosis af
C0004238|000|rheumatic af
C0004238|000|chf with af
C0004238|000|hfpef with af
C0004238|000|hfref with af
C0004238|000|chf/af
C0004238|000|hf/af
C0004238|000|dilated cardiomyopathy with af
C0004238|000|dcm/af
C0004238|000|cardioembolic af
C0004238|000|thromboembolic af
C0004238|000|thyrotoxic af
C0004238|000|hyperthyroid af
C0004238|000|thyrotoxic atrial fibrillation
C0004238|000|post-cardiac surgery af
C0004238|000|surgery-induced af
C0004238|000|postablation af
C0004238|000|post-ablation a-fib
C0004238|000|lone af
C0004238|000|cryptogenic af
C0004238|000|familial af
C0004238|000|inherited af
C0004238|000|idiopathic af
C0004238|000|spontaneous af
C0004238|000|secondary to sepsis af
C0004238|000|sepsis-associated af
C0004238|000|post-mi af
C0004238|000|post infarct af
C0004238|000|post cabg af
C0004238|000|cabg-related af
C0004238|000|post-op a-fib
C0004238|000|perioperative af
C0004238|000|renal failure with af
C0004238|000|af in ckd
C0004238|000|esrd with af
C0004238|000|dialysis-associated af
C0004238|000|copd-related af
C0004238|000|obstructive sleep apnea with af
C0004238|000|osa with af
C0004238|000|af in elderly
C0004238|000|degenerative af
C0004238|000|afiv
C0004238|000|a fib
C0004238|000|afib episode
C0004238|000|asx af
C0004238|000|parox af
C0004238|000|sym af
C0004238|000|asymp af
C0004238|000|atrial fib episode
C0004238|000|beta-blocker controlled af
C0004238|000|rate-controlled af
C0004238|000|rhythm-controlled af
C0004238|000|af on anticoagulation
C0004238|000|af on oac
C0004238|000|af with stroke
C0004238|000|af with embolism
C0004238|000|embolic a-fib
C0004238|000|af of unknown cause
C0004238|000|af post anaesthesia
C0004238|000|af on ecg
C0004238|000|ecg: af
C0004238|000|telemetry: af
C0004238|000|holter: af
C0004238|000|atrial fib rvr
C0004238|000|fib w/ rvr
C0004238|000|af/svr
C0004238|000|tachy af
C0004238|000|persistent afib
C0004238|000|chronic afib
C0004238|000|recurring afib
C0004238|000|long-term afib
C0004238|000|persistent a fib
C0004238|000|intermittent af
C0004238|000|episodes of af
C0004238|000|brief af
C0004238|000|asx atrial fib
C0004238|000|supraventricular af
C0015672|000|fatigue
C0015672|000|fatigued
C0015672|000|fatiging
C0015672|000|fatigability
C0015672|000|easy fatigability
C0015672|000|early fatigability
C0015672|000|increased fatigability
C0015672|000|severe fatigue
C0015672|000|chronic fatigue
C0015672|000|malaise
C0015672|000|lassitude
C0015672|000|tired
C0015672|000|tiredness
C0015672|000|easily tired
C0015672|000|exercise intolerance
C0015672|000|dec exercise tolerance
C0015672|000|poor exercise tolerance
C0015672|000|exertional fatigue
C0015672|000|exercise-induced fatigue
C0015672|000|post-exertional fatigue
C0015672|000|weakness
C0015672|000|generalized weakness
C0015672|000|muscle weakness
C0015672|000|subjective weakness
C0015672|000|lethargy
C0015672|000|lethargic
C0015672|000|exhaustion
C0015672|000|exhausted
C0015672|000|low energy
C0015672|000|decreased energy
C0015672|000|dec energy
C0015672|000|loss of energy
C0015672|000|easy exhaustion
C0015672|000|quickly exhausted
C0015672|000|no stamina
C0015672|000|reduced stamina
C0015672|000|low stamina
C0015672|000|weariness
C0015672|000|worn out
C0015672|000|drained
C0015672|000|sluggishness
C0015672|000|sluggish
C0015672|000|slowness
C0015672|000|nonrestorative sleep
C0015672|000|non-restful sleep
C0015672|000|daytime sleepiness
C0015672|000|somnolence
C0015672|000|drowsiness
C0015672|000|sleepiness
C0015672|000|poor tolerance to activity
C0015672|000|activity intolerance
C0015672|000|easy fatigued
C0015672|000|subjective fatigue
C0015672|000|chemo-induced fatigue
C0015672|000|chemotherapy-related fatigue
C0015672|000|ca fatigue
C0015672|000|post-chemo fatigue
C0015672|000|crf
C0015672|000|cancer fatigue
C0015672|000|radiation-induced fatigue
C0015672|000|anemia-associated fatigue
C0015672|000|anemic fatigue
C0015672|000|hf fatigue
C0015672|000|chf fatigue
C0015672|000|heart failure fatigue
C0015672|000|ischemic fatigue
C0015672|000|low cardiac output fatigue
C0015672|000|amyloid fatigue
C0015672|000|amyloidosis-related fatigue
C0015672|000|valvular fatigue
C0015672|000|hypertensive fatigue
C0015672|000|htn fatigue
C0015672|000|htn-related fatigue
C0015672|000|myocarditis fatigue
C0015672|000|tachycardia-induced fatigue
C0015672|000|arrhythmia-related fatigue
C0015672|000|postviral fatigue
C0015672|000|viral fatigue
C0015672|000|infectious fatigue
C0015672|000|post-covid fatigue
C0015672|000|covid fatigue
C0015672|000|me/cfs
C0015672|000|chronic fatigue syndrome
C0015672|000|post-infectious fatigue
C0015672|000|hiv-related fatigue
C0015672|000|apls fatigue
C0015672|000|ppcm fatigue
C0015672|000|peripartum fatigue
C0015672|000|pregnancy-induced fatigue
C0015672|000|postpartum fatigue
C0015672|000|endocrine fatigue
C0015672|000|thyroid-related fatigue
C0015672|000|hypothyroid fatigue
C0015672|000|hypothyroidism fatigue
C0015672|000|adrenal fatigue
C0015672|000|addison’s fatigue
C0015672|000|diabetic fatigue
C0015672|000|renal fatigue
C0015672|000|ckd fatigue
C0015672|000|renal failure fatigue
C0015672|000|hepatic fatigue
C0015672|000|liver failure fatigue
C0015672|000|cld fatigue
C0015672|000|malignancy fatigue
C0015672|000|sle fatigue
C0015672|000|ra fatigue
C0015672|000|ms fatigue
C0015672|000|neuromuscular fatigue
C0015672|000|depression-related fatigue
C0015672|000|psychogenic fatigue
C0015672|000|mental fatigue
C0015672|000|cognitive fatigue
C0015672|000|fibromyalgia fatigue
C0015672|000|pain-related fatigue
C0015672|000|post-concussion fatigue
C0015672|000|tbi fatigue
C0015672|000|chronic disease fatigue
C0015672|000|post-surgical fatigue
C0015672|000|post-op fatigue
C0015672|000|drug-induced fatigue
C0015672|000|medication-related fatigue
C0015672|000|antidepressant fatigue
C0015672|000|antipsychotic fatigue
C0015672|000|sleep apnea fatigue
C0015672|000|osa fatigue
C0015672|000|csa fatigue
C0015672|000|night sweats and fatigue
C0015672|000|migrainous fatigue
C0015672|000|fatigue of unknown etiology
C0015672|000|idiopathic fatigue
C0015672|000|ebv fatigue
C0015672|000|lyme fatigue
C0015672|000|rheumatologic fatigue
C0015672|000|crps fatigue
C0015672|000|copd fatigue
C0015672|000|pulmonary fatigue
C0015672|000|respiratory fatigue
C0015672|000|disease-related fatigue
C0015672|000|tired out
C0015672|000|wiped out
C0015672|000|run down
C0015672|000|flagging
C0015672|000|lack of pep
C0015672|000|lack of vigor
C0015672|000|slowed down
C0015672|000|lacks energy
C0015672|000|needs naps
C0015672|000|falls asleep during day
C0015672|000|reduced activity tolerance
C0015672|000|reduced functional capacity
C0015672|000|cannot keep up usual activity
C0015672|000|mental exhaustion
C0015672|000|physical exhaustion
C0015672|000|overwhelming fatigue
C0015672|000|burnout
C0015672|000|asthenia
C0015672|000|listlessness
C0015672|000|debilitation
C0015672|000|debilitated
C0015672|000|profound fatigue
C0015672|000|significant fatigue
C0015672|000|marked fatigue
C0015672|000|extreme fatigue
C0015672|000|incapacitating fatigue
C0015672|000|insufficient energy
C0015672|000|difficulty completing tasks
C0015672|000|reports fatigue
C0015672|000|pt c/o fatigue
C0015672|000|c/o tiredness
C0015672|000|sensation of weakness
C0015672|000|decreased activity
C0015672|000|cannot finish adls
C0015672|000|decreased job performance
C0015672|000|not feeling rested
C0015672|000|persistent tiredness
C0015672|000|ongoing fatigue
C0015672|000|constant fatigue
C0015672|000|intermittent fatigue
C0015672|000|periodic fatigue
C0015672|000|worsening fatigue
C0015672|000|recurrent fatigue
C0015672|000|energy deficit
C0015672|000|vitality loss
C0015672|000|weakness
C0015672|000|generalized weakness
C0015672|000|focal weakness
C0015672|000|muscle weakness
C0015672|000|proximal weakness
C0015672|000|distal weakness
C0015672|000|asthenia
C0015672|000|paresis
C0015672|000|hemiparesis
C0015672|000|paraparesis
C0015672|000|quadriparesis
C0015672|000|tetraparesis
C0015672|000|myopathy
C0015672|000|fatigue
C0015672|000|malaise
C0015672|000|decreased strength
C0015672|000|low strength
C0015672|000|diminished strength
C0015672|000|loss of strength
C0015672|000|power loss
C0015672|000|reduced power
C0015672|000|motor deficit
C0015672|000|motor impairment
C0015672|000|flaccidity
C0015672|000|flaccid muscles
C0015672|000|muscular fatigue
C0015672|000|exertional fatigue
C0015672|000|neuromuscular weakness
C0015672|000|hyposthenia
C0015672|000|nm weakness
C0015672|000|decreased grip strength
C0015672|000|sluggish muscle response
C0015672|000|muscle atony
C0015672|000|muscle hypotonia
C0015672|000|floppy muscles
C0015672|000|muscle insufficiency
C0015672|000|myasthenia
C0015672|000|ppcm-related weakness
C0015672|000|cva-related weakness
C0015672|000|stroke-related weakness
C0015672|000|ischemic weakness
C0015672|000|nonischemic weakness
C0015672|000|chemo-induced weakness
C0015672|000|drug-induced weakness
C0015672|000|myocarditis-related weakness
C0015672|000|valvular-related weakness
C0015672|000|hypertensive weakness
C0015672|000|amyloid weakness
C0015672|000|tachycardia-induced weakness
C0015672|000|als-related weakness
C0015672|000|ms-related weakness
C0015672|000|parkinsonian weakness
C0015672|000|alcoholic weakness
C0015672|000|critical illness weakness
C0015672|000|periodic paralysis
C0015672|000|central weakness
C0015672|000|peripheral weakness
C0015672|000|monoparesis
C0015672|000|paresis rle
C0015672|000|paresis lle
C0015672|000|paresis rue
C0015672|000|paresis lue
C0015672|000|le weakness
C0015672|000|rle weakness
C0015672|000|lle weakness
C0015672|000|ue weakness
C0015672|000|rue weakness
C0015672|000|lue weakness
C0015672|000|diffuse weakness
C0015672|000|bilateral weakness
C0015672|000|unilateral weakness
C0015672|000|r-sided weakness
C0015672|000|l-sided weakness
C0015672|000|impaired muscle strength
C0015672|000|mobility impairment
C0015672|000|ambulatory weakness
C0015672|000|transient weakness
C0015672|000|chronic weakness
C0015672|000|acute weakness
C0015672|000|subjective weakness
C0015672|000|objective weakness
C0015672|000|myotonia
C0015672|000|em weakness
C0015672|000|functional weakness
C0015672|000|secondary weakness
C0015672|000|progressive weakness
C0015672|000|persistent weakness
C0015672|000|episodic weakness
C0015672|000|muscle deficit
C0015672|000|neuropathic weakness
C0015672|000|myopathic weakness
C0015672|000|limb weakness
C0015672|000|down-going strength
C0015672|000|paresis limb
C0015672|000|paresis extremity
C0015672|000|motor weakness
C0015672|000|loss of muscle function
C0015672|000|muscle deterioration
C0015672|000|muscle debility
C0015672|000|muscle flaccidity
C0015672|000|gait weakness
C0015672|000|muscle sluggishness
C0015672|000|frank weakness
C0015672|000|mild weakness
C0015672|000|moderate weakness
C0015672|000|marked weakness
C0015672|000|severe weakness
C0015672|000|pml-related weakness
C0015672|000|gbs-related weakness
C0015672|000|mnd weakness
C0015672|000|cidp-related weakness
C0015672|000|inflammatory weakness
C0015672|000|immune-mediated weakness
C0015672|000|cachectic weakness
C0015672|000|paraneoplastic weakness
C0015672|000|disuse weakness
C0015672|000|immobility-related weakness
C0015672|000|respiratory muscle weakness
C0015672|000|oculomotor weakness
C0015672|000|bulbar weakness
C0015672|000|facial weakness
C0015672|000|cranial nerve weakness
C0015672|000|truncal weakness
C0015672|000|core weakness
C0015672|000|hand weakness
C0015672|000|wrist drop
C0015672|000|foot drop
C0015672|000|muscle fatigability
C0015672|000|easy fatigability
C0015672|000|pem (post-exertional malaise)
C0015672|000|floppy baby
C0015672|000|motor neuron weakness
C0015672|000|neurogenic weakness
C0015672|000|recurrent weakness
C0015672|000|fluctuant weakness
C0015672|000|waxing/waning weakness
C0015672|000|emg-documented weakness
C0015672|000|exercise-induced weakness
C0015672|000|overuse weakness
C0015672|000|debilitation
C0015672|000|muscular debility
C0015672|000|myasthenic symptoms
C0015672|000|hypotonicity
C0015672|000|decreased tone
C0015672|000|drop attacks
C0015672|000|loss muscle bulk
C0015672|000|atrophic weakness
C0015672|000|lateralizing weakness
C0015672|000|symmetric weakness
C0015672|000|asymmetric weakness
C0015672|000|spastic weakness
C0015672|000|nonspastic weakness
C0015672|000|limb drift
C0015672|000|pronator drift
C0015672|000|clumsiness
C0015672|000|unsteady
C0015672|000|loss of antigravity strength
C0015672|000|muscle impairment
C0015672|000|poor muscle performance
C0015672|000|impaired performance
C0015672|000|decline muscle strength
C0015672|000|mechanical weakness
C0015672|000|myotoxicity
C0015672|000|toxic myopathy
C0015672|000|steroid-induced weakness
C0015672|000|corticosteroid myopathy
C0015672|000|paraplegic weakness
C0015672|000|plegic weakness
C0015672|000|flaccid paresis
C0015672|000|hypotonic weakness
C0015672|000|lower limb weakness
C0015672|000|upper limb weakness
C0015672|000|speech weakness
C0015672|000|dysarthric weakness
C0015672|000|pharyngeal weakness
C0015672|000|lingual weakness
C0015672|000|tongue weakness
C0015672|000|neck flexion weakness
C0015672|000|neck extension weakness
C0015672|000|axial weakness
C0015672|000|presynaptic weakness
C0015672|000|postsynaptic weakness
C0015672|000|distal limb weakness
C0015672|000|proximal limb weakness
C0015672|000|hand grip weakness
C0015672|000|paresis ues
C0015672|000|paresis les
C0015672|000|progressive myopathy
C0015672|000|myopathy nos
C0015672|000|myositis-related weakness
C0015672|000|limb heaviness
C0015672|000|heavy limbs
C0015672|000|muscle heaviness
C0015672|000|floppy infant
C0015672|000|myasthenic weakness
C0015672|000|neoplasm-related weakness
C0015672|000|critical illness myopathy
C0015672|000|systemic weakness
C0015672|000|pandysautonomia weakness
C5543391|000|low appetite
C5543391|000|↓ appetite
C5543391|000|decreased appetite
C5543391|000|dec appetite
C5543391|000|↓ po intake
C5543391|000|po intake ↓
C5543391|000|poor appetite
C5543391|000|reduced appetite
C5543391|000|loss of appetite
C5543391|000|appetite loss
C5543391|000|appetite ↓
C5543391|000|no appetite
C5543391|000|anorexia
C5543391|000|anorexic
C5543391|000|anorexia nervosa
C5543391|000|poor oral intake
C5543391|000|↓ oral intake
C5543391|000|low oral intake
C5543391|000|oral intake ↓
C5543391|000|diminished appetite
C5543391|000|diminished po intake
C5543391|000|appetite off
C5543391|000|avoiding food
C5543391|000|not eating well
C5543391|000|not eating
C5543391|000|decreased eating
C5543391|000|eating less
C5543391|000|appetite suppression
C5543391|000|anorexia (chemo-induced)
C5543391|000|chemo-induced anorexia
C5543391|000|chemo-induced appetite loss
C5543391|000|loss of appetite (chemo)
C5543391|000|appetite change
C5543391|000|poor po
C5543391|000|↓ po
C5543391|000|po poor
C5543391|000|s/p chemo ↓ appetite
C5543391|000|appetite poor
C5543391|000|low caloric intake
C5543391|000|↓ caloric intake
C5543391|000|hyporexia
C5543391|000|hyporexic
C5543391|000|poor feeding
C5543391|000|reduced feeding
C5543391|000|failure to thrive (ftt)
C5543391|000|ftt
C5543391|000|cachexia
C5543391|000|cancer cachexia
C5543391|000|tumor-induced anorexia
C5543391|000|nonischemic anorexia
C5543391|000|ischemic anorexia
C5543391|000|anorexia (myocarditis)
C5543391|000|tachycardia-induced anorexia
C5543391|000|myocarditis-related poor appetite
C5543391|000|chf-related loss of appetite
C5543391|000|valvular disease ↓ appetite
C5543391|000|appetite down
C5543391|000|poor intake
C5543391|000|decreased intake
C5543391|000|npo except meds
C5543391|000|intake less than baseline
C5543391|000|low nutritional intake
C5543391|000|food aversion
C5543391|000|feeding aversion
C5543391|000|reduced nutritional intake
C5543391|000|↓ interest in food
C5543391|000|reluctant to eat
C5543391|000|not hungry
C5543391|000|inappetent
C5543391|000|appetite suppressed
C5543391|000|self-restricted dietary intake
C5543391|000|poor nutrition
C5543391|000|voluntary starvation
C5543391|000|intentional anorexia
C5543391|000|starvation (anorexia)
C5543391|000|poor intake (ppcm)
C5543391|000|amyloidosis-related appetite loss
C5543391|000|amyloidosis poor appetite
C5543391|000|inadequate po intake
C5543391|000|low po
C5543391|000|low food consumption
C5543391|000|eating < normal
C5543391|000|intake < normal
C5543391|000|↓ food consumption
C5543391|000|diminished desire to eat
C5543391|000|unable to tolerate po
C5543391|000|appetite lacking
C5543391|000|decreased desire for food
C5543391|000|loss of interest in eating
C5543391|000|skipping meals
C5543391|000|refusing meals
C5543391|000|using appetite suppressants
C5543391|000|gi-related ↓ appetite
C5543391|000|hepatic anorexia
C5543391|000|heart failure anorexia
C5543391|000|cardiac cachexia
C5543391|000|ckd-related anorexia
C5543391|000|esrd-related poor appetite
C5543391|000|dialysis-related ↓ appetite
C5543391|000|uremic anorexia
C5543391|000|copd-related ↓ appetite
C5543391|000|hiv-related anorexia
C5543391|000|infection-related loss of appetite
C5543391|000|sepsis anorexia
C5543391|000|tb-related poor appetite
C5543391|000|anorexia secondary to disease
C5543391|000|malignancy-related ↓ appetite
C5543391|000|oncologic anorexia
C5543391|000|appetite complaint
C5543391|000|reduced caloric intake
C5543391|000|nutrition intake suboptimal
C5543391|000|nutrition: poor
C5543391|000|nutrition: decreased
C5543391|000|eats very little
C5543391|000|minimal po intake
C5543391|000|↓ consumption
C5543391|000|low dietary intake
C5543391|000|dietary intake reduced
C5543391|000|unable to eat
C5543391|000|feeding difficulty
C5543391|000|reluctance to feed
C5543391|000|anorexia (psychiatric)
C5543391|000|geriatric anorexia
C5543391|000|pediatric poor feeding
C5543391|000|hunger absent
C5543391|000|non-volitional ↓ intake
C5543391|000|self-limited po
C5543391|000|voluntarily not eating
C5543391|000|hypophagia
C5543391|000|hypophagic
C5543391|000|prn appetite loss
C5543391|000|drug-induced anorexia
C5543391|000|opioid-induced ↓ appetite
C5543391|000|antibiotic-induced ↓ appetite
C5543391|000|ssris - appetite loss
C5543391|000|steroid-induced ↓ appetite
C5543391|000|appetite suppressed (rx)
C5543391|000|stress-induced anorexia
C5543391|000|depression-related decreased appetite
C5543391|000|anxiety-related anorexia
C5543391|000|po intolerance
C5543391|000|unable to tolerate oral intake
C5543391|000|failure to eat
C5543391|000|refusal to eat
C5543391|000|appetite reduced
C5543391|000|appetite significantly ↓
C5543391|000|sarcopenia-related poor intake
C5543391|000|impaired appetite
C5543391|000|low feeding drive
C5543391|000|early satiety
C5543391|000|no desire for food
C5543391|000|satiety at low volumes
C5543391|000|perceived anorexia
C5543391|000|progressive decrease in appetite
C5543391|000|acute onset anorexia
C5543391|000|chronic poor appetite
C5543391|000|recurrent anorexia
C5543391|000|appetite disturbance
C5543391|000|low interest in food
C5543391|000|gastrointestinal symptoms - poor appetite
C5543391|000|post-op ↓ appetite
C5543391|000|post-infectious anorexia
C5543391|000|postpartum poor appetite
C5543391|000|pregnancy-related appetite loss
C5543391|000|appetite off since illness
C5543391|000|withdrew from eating
C5543391|000|low po tolerance
C5543391|000|poor caloric intake
C5543391|000|appetite not present
C5543391|000|cannot tolerate diet
C5543391|000|appetite declining
C5543391|000|eating reluctance
C5543391|000|no feeding
C5543391|000|neglecting meals
C5543391|000|adhf-related ↓ appetite
C5543391|000|low po desire
C5543391|000|lack of hunger
C5543391|000|reduced food preference
C5543391|000|reduced desire for food
C0003123|000|anorexia
C0003123|000|anorexic
C0003123|000|↓ appetite
C0003123|000|decreased appetite
C0003123|000|loss of appetite
C0003123|000|poor appetite
C0003123|000|reduced appetite
C0003123|000|anorexia nervosa
C0003123|000|cancer anorexia
C0003123|000|chemo-induced anorexia
C0003123|000|drug-induced anorexia
C0003123|000|appetite loss
C0003123|000|appetite suppression
C0003123|000|no appetite
C0003123|000|failure to eat
C0003123|000|refusing food
C0003123|000|not eating
C0003123|000|appetite reduction
C0003123|000|inappetence
C0003123|000|hyporexia
C0003123|000|appetite decline
C0003123|000|diminished appetite
C0003123|000|lack of appetite
C0003123|000|poor po intake
C0003123|000|anorexia-cachexia
C0003123|000|a/n
C0003123|000|a/nv
C0003123|000|chf-related anorexia
C0003123|000|ckd-related anorexia
C0003123|000|esrd anorexia
C0003123|000|uremic anorexia
C0003123|000|gi-induced anorexia
C0003123|000|infectious anorexia
C0003123|000|psychogenic anorexia
C0003123|000|depression-related anorexia
C0003123|000|hepatic anorexia
C0003123|000|liver disease anorexia
C0003123|000|dementia anorexia
C0003123|000|dementia-related decreased appetite
C0003123|000|appetite off
C0003123|000|not interested in food
C0003123|000|patient not eating
C0003123|000|voluntary food restriction
C0003123|000|starvation
C0003123|000|no po
C0003123|000|↓ oral intake
C0003123|000|not tolerating po
C0003123|000|↓ food intake
C0003123|000|minimal intake
C0003123|000|reduced po intake
C0003123|000|decreased po
C0003123|000|refusal to eat
C0575081|000|gait abnormality
C0575081|000|abnormal gait
C0575081|000|gait disturbance
C0575081|000|abnormal gait pattern
C0575081|000|disordered gait
C0575081|000|ataxic gait
C0575081|000|gait ataxia
C0575081|000|unsteady gait
C0575081|000|walking difficulty
C0575081|000|disturbed ambulation
C0575081|000|abnormal ambulation
C0575081|000|ambulatory dysfunction
C0575081|000|abnormal walking
C0575081|000|impaired gait
C0575081|000|gait impairment
C0575081|000|ambulatory impairment
C0575081|000|difficulty walking
C0575081|000|impaired ambulation
C0575081|000|abnormal locomotion
C0575081|000|locomotor abnormality
C0575081|000|gait instability
C0575081|000|instability walking
C0575081|000|unstable gait
C0575081|000|gait dyspraxia
C0575081|000|shuffling gait
C0575081|000|festinating gait
C0575081|000|parkinsonian gait
C0575081|000|spastic gait
C0575081|000|spastic-ataxic gait
C0575081|000|hemiplegic gait
C0575081|000|hemiparetic gait
C0575081|000|diplegic gait
C0575081|000|scissoring gait
C0575081|000|scissor gait
C0575081|000|trendelenburg gait
C0575081|000|waddling gait
C0575081|000|cerebellar gait
C0575081|000|sensory ataxia
C0575081|000|apraxic gait
C0575081|000|myopathic gait
C0575081|000|steppage gait
C0575081|000|neuropathic gait
C0575081|000|foot drop gait
C0575081|000|paraparetic gait
C0575081|000|high-stepping gait
C0575081|000|magnetic gait
C0575081|000|hypokinetic gait
C0575081|000|bradykinetic gait
C0575081|000|tabetic gait
C0575081|000|choreiform gait
C0575081|000|antalgic gait
C0575081|000|limping gait
C0575081|000|limp
C0575081|000|walking abnormality
C0575081|000|walking disturbance
C0575081|000|abnl gait
C0575081|000|gait abnl
C0575081|000|gait dis
C0575081|000|gait dist
C0575081|000|impaired walking
C0575081|000|mobility impairment
C0575081|000|mobility abnormality
C0575081|000|decreased mobility
C0575081|000|gait dysfunction
C0575081|000|gait unsteadiness
C0575081|000|wide-based gait
C0575081|000|narrow-based gait
C0575081|000|small steps gait
C0575081|000|short stride gait
C0575081|000|gait freezing
C0575081|000|gait block
C0575081|000|propulsive gait
C0575081|000|paretic gait
C0575081|000|staggering gait
C0575081|000|drunken gait
C0575081|000|elderly gait disturbance
C0575081|000|frontal gait disorder
C0575081|000|gait disorder nos
C0575081|000|abnormal gait nos
C0575081|000|gait disturbance nos
C0575081|000|difficulty ambulating
C0575081|000|impaired gross mobility
C0575081|000|slow gait
C0575081|000|slowness walking
C0575081|000|gait slowness
C0575081|000|cautious gait
C0575081|000|gait hesitation
C0575081|000|equinus gait
C0575081|000|toe-walking
C0575081|000|toe gait
C0575081|000|calcaneal gait
C0575081|000|heel-walking
C0575081|000|clumsy gait
C0575081|000|abnl ambulation
C0575081|000|ms-related gait dysfunction
C0575081|000|parkinson's gait
C0575081|000|hemiplegic walking
C0575081|000|functional gait disorder
C0575081|000|conversion gait
C0575081|000|psychogenic gait
C0575081|000|malingered gait
C0575081|000|tremor during gait
C0575081|000|dystonic gait
C0575081|000|spastic-hemiplegic gait
C0575081|000|flaccid gait
C0575081|000|choreaform gait
C0575081|000|basal ganglia gait disorder
C0575081|000|extrapyramidal gait disorder
C0575081|000|gait apraxia
C0575081|000|gait difficulty
C0575081|000|abnormal stride
C0575081|000|gait deviation
C0575081|000|gait change
C0575081|000|gait deficit
C0575081|000|poor gait
C0575081|000|altered gait
C0575081|000|altered ambulation
C0575081|000|disrupted gait
C0575081|000|gait impairment due to stroke
C0575081|000|post-stroke gait
C0575081|000|ischemic gait abnormality
C0575081|000|chemo-induced gait abnormality
C0575081|000|myelopathy-related gait disorder
C0575081|000|radiculopathy gait abnormality
C0575081|000|als-related gait abnormality
C0575081|000|motor neuron gait deficit
C0575081|000|pyramidal gait
C0575081|000|spinal gait disturbance
C0575081|000|cerebral palsy gait
C0575081|000|cp gait
C0575081|000|demyelinating gait
C0575081|000|peripheral neuropathy gait
C0575081|000|diabetic gait disturbance
C0575081|000|amyloid gait abnormality
C0575081|000|hypertensive gait disorder
C0575081|000|valvular gait disorder
C0575081|000|tachycardia-induced gait abnormality
C0575081|000|ppcm gait abnormality
C0575081|000|myocarditis gait abnormality
C0575081|000|mixed pattern gait
C0575081|000|sensory-motor gait disturbance
C0575081|000|posterior column gait disorder
C0575081|000|spastic-paraparetic gait
C0575081|000|bilateral gait disturbance
C0575081|000|bilateral leg gait abnormality
C0575081|000|spastic quadriparetic gait
C0575081|000|quadriparetic gait
C0575081|000|unmotivated gait
C0575081|000|weak gait
C0575081|000|loss of gait automation
C0575081|000|frontal ataxia
C0575081|000|subcortical gait disturbance
C0575081|000|akinetic gait
C0575081|000|hypometric gait
C0575081|000|dyskinetic gait
C0575081|000|hyperkinetic gait
C0575081|000|swaying gait
C0575081|000|leaning gait
C0575081|000|lateralized gait
C0575081|000|ill-compensated gait
C0575081|000|postural gait abnormality
C0575081|000|drop foot gait
C0575081|000|hemiparetic walking
C0575081|000|toe drag gait
C0575081|000|step-page gait
C0575081|000|stooped gait
C0575081|000|stiff-legged gait
C0575081|000|genu recurvatum gait
C0575081|000|myotonic gait
C0575081|000|ataxia
C0575081|000|gmf dysfunction
C0575081|000|gmf deficit
C0575081|000|trendelenburg sign
C0575081|000|incoordinated gait
C0575081|000|nonphysiologic gait
C0575081|000|friction gait
C0575081|000|gait deviation due to spasticity
C0575081|000|spasticity-related gait change
C0575081|000|spastic diplegic gait
C0575081|000|dysfunctional stride
C0575081|000|gait variance
C0241981|000|impaired balance
C0241981|000|balance impairment
C0241981|000|unsteady gait
C0241981|000|gait instability
C0241981|000|ataxia
C0241981|000|vestibular dysfunction
C0241981|000|loss of balance
C0241981|000|postural instability
C0241981|000|impaired coordination
C0241981|000|equilibrium disturbance
C0241981|000|gait disturbance
C0241981|000|unsteadiness
C0241981|000|dizziness
C0241981|000|disequilibrium
C0241981|000|vertigo
C0241981|000|unsteady on feet
C0241981|000|wobbling gait
C0241981|000|staggering
C0241981|000|romberg positive
C0241981|000|wide-based gait
C0241981|000|abnormal gait
C0241981|000|waddling gait
C0241981|000|lurching gait
C0241981|000|drunken gait
C0241981|000|gait ataxia
C0241981|000|impaired proprioception
C0241981|000|impaired vestibular function
C0241981|000|labyrinthine dysfunction
C0241981|000|cerebellar ataxia
C0241981|000|sensory ataxia
C0241981|000|vestibular ataxia
C0241981|000|spinocerebellar ataxia
C0241981|000|paraparesis
C0241981|000|spastic gait
C0241981|000|toe-walking
C0241981|000|impairment of equilibrium
C0241981|000|impaired stance
C0241981|000|swaying
C0241981|000|gait abnormality
C0241981|000|shuffling gait
C0241981|000|parkinsonian gait
C0241981|000|gait deviation
C0241981|000|sway-positive
C0241981|000|antalgic gait
C0241981|000|hemiparetic gait
C0241981|000|ataxic gait
C0241981|000|impaired ambulation
C0241981|000|poor balance
C0241981|000|abnormal tandem gait
C0241981|000|abnormal heel-to-toe walk
C0241981|000|impaired tandem gait
C0241981|000|instability
C0241981|000|gait disorder
C0241981|000|gait unsteadiness
C0241981|000|marching unsteadily
C0241981|000|perceived imbalance
C0241981|000|oscillopsia
C0241981|000|feelings of imbalance
C0241981|000|impaired postural control
C0241981|000|abnormal posture
C0241981|000|bilateral leg unsteadiness
C0241981|000|loss of proprioception
C0241981|000|falling tendencies
C0241981|000|near falls
C0241981|000|off-balance
C0241981|000|loss of stability
C0241981|000|gait uncoordination
C0241981|000|drifting to side
C0241981|000|proprioceptive deficit
C0241981|000|sway on standing
C0241981|000|impaired romberg
C0241981|000|positive romberg
C0241981|000|disordered equilibrium
C0241981|000|gait dyspraxia
C0241981|000|dysmetria
C0241981|000|dysequilibrium
C0241981|000|locomotor ataxia
C0241981|000|veering
C0241981|000|poor righting reflex
C0241981|000|abnormal righting response
C0241981|000|truncal ataxia
C0241981|000|hypotonic gait
C0241981|000|gait freezing
C0241981|000|festination
C0241981|000|drop attacks
C0241981|000|frequent stumbles
C0241981|000|frequent falls
C0241981|000|abnormal gait mechanics
C0241981|000|limb incoordination
C0241981|000|balance deficit
C0241981|000|balance disorder
C0241981|000|compromised balance
C0241981|000|equilibrium disorder
C0241981|000|abnormal balance
C0241981|000|impaired verticality
C0241981|000|standing instability
C0241981|000|abnormal balance test
C0241981|000|proprioceptive gait disorder
C0241981|000|myopathy gait
C0241981|000|neuropathic gait
C0241981|000|steppage gait
C0241981|000|acute vestibulopathy
C0241981|000|central vestibulopathy
C0241981|000|peripheral vestibulopathy
C0241981|000|cerebellopathy
C0241981|000|ischemic ataxia
C0241981|000|nonischemic ataxia
C0241981|000|stroke-related instability
C0241981|000|tbi-related balance loss
C0241981|000|cva with gait disturbance
C0241981|000|ms-related ataxia
C0241981|000|parkinson’s gait disturbance
C0241981|000|chemo-induced ataxia
C0241981|000|medication-induced imbalance
C0241981|000|alcohol-induced ataxia
C0241981|000|diabetic ataxia
C0241981|000|amyloid neuropathy gait
C0241981|000|thiamine-deficient ataxia
C0241981|000|vitamin b12 deficiency gait
C0241981|000|myelopathy-induced gait impairment
C0241981|000|spinal stenosis–related balance loss
C0241981|000|peripheral neuropathy–related imbalance
C0241981|000|sensory neuropathy gait
C0241981|000|tachycardia-induced syncope with falls
C0241981|000|ppcm-related unsteady gait
C0241981|000|chf with instability
C0241981|000|hypertensive encephalopathy ataxia
C0241981|000|cerebellar infarct with imbalance
C0241981|000|vertebrobasilar insufficiency with ataxia
C0241981|000|valvular disease with falls
C0241981|000|meniere’s disease imbalance
C0241981|000|bppv imbalance
C0241981|000|ototoxicity with gait disturbance
C0241981|000|presbystasis
C0241981|000|areflexia with unsteady gait
C0241981|000|ortho hypotension with falls
C0241981|000|acute labyrinthitis
C0241981|000|chronic imbalance
C0241981|000|idiopathic ataxia
C0241981|000|post-ictal unsteadiness
C0241981|000|post-surgical imbalance
C0241981|000|age-related imbalance
C0241981|000|impaired walk
C0241981|000|coordination deficit
C0241981|000|uncoordinated gait
C0241981|000|disordered gait
C0241981|000|impaired locomotion
C0241981|000|impaired walking stability
C0241981|000|tripping easily
C0241981|000|impaired stance control
C0241981|000|marked gait disturbance
C0241981|000|walks with assistance
C0241981|000|requires mobility aid
C0241981|000|frequent wall walking
C0241981|000|unstable gait
C0241981|000|instability on ambulation
C0241981|000|poor postural stability
C0241981|000|unsteady when turning
C0241981|000|unsteady standing
C0241981|000|poor dynamic balance
C0241981|000|deficient balance response
C0241981|000|impaired dynamic equilibrium
C0241981|000|imbalance
C0241981|000|bos-wide gait
C0241981|000|need for assistive device due to balance
C0241981|000|use of cane for balance
C1405979|000|radiation necrosis
C1405979|000|radiation-induced necrosis
C1405979|000|post-radiation necrosis
C1405979|000|postirradiation necrosis
C1405979|000|radionecrosis
C1405979|000|radiation-related necrosis
C1405979|000|rn
C1405979|000|rt necrosis
C1405979|000|radio-necrosis
C1405979|000|irradiation necrosis
C1405979|000|necrosis secondary to radiation
C1405979|000|necrosis d/t radiation
C1405979|000|necrosis s/p radiation
C1405979|000|necrosis d/t rt
C1405979|000|necrosis s/p rt
C1405979|000|necrosis s/p irradiation
C1405979|000|post-radiotherapy necrosis
C1405979|000|radiotherapy necrosis
C1405979|000|necrosis following ionizing radiation
C1405979|000|ionizing radiation necrosis
C1405979|000|necrosis due to radiotherapy
C1405979|000|post-rt necrosis
C1405979|000|radiation necrotic changes
C1405979|000|radionecrotic lesion
C1405979|000|radiation injury with necrosis
C1405979|000|radiation effect necrosis
C1405979|000|secondary radiation necrosis
C1405979|000|delayed radiation necrosis
C1405979|000|delayed radionecrosis
C1405979|000|late rt necrosis
C1405979|000|late radiation necrosis
C1405979|000|chronic radiation necrosis
C1405979|000|chronic radionecrosis
C1405979|000|focal radiation necrosis
C1405979|000|multifocal radiation necrosis
C1405979|000|gliocentric radiation necrosis
C1405979|000|nonischemic radiation necrosis
C1405979|000|ischemic radiation necrosis
C1405979|000|necrosis due to therapeutic irradiation
C1405979|000|therapy-induced necrosis
C1405979|000|treatment-induced necrosis
C1405979|000|necrosis post-external beam rt
C1405979|000|necrosis secondary to ebrt
C1405979|000|ebrt necrosis
C1405979|000|gamma knife necrosis
C1405979|000|stereotactic radiosurgery necrosis
C1405979|000|srs necrosis
C1405979|000|srt necrosis
C1405979|000|sbrt necrosis
C1405979|000|cns radiation necrosis
C1405979|000|brain radiation necrosis
C1405979|000|cerebral radiation necrosis
C1405979|000|myocardial radiation necrosis
C1405979|000|hepatic radiation necrosis
C1405979|000|pancreatic radiation necrosis
C1405979|000|soft tissue radiation necrosis
C1405979|000|cutaneous radiation necrosis
C1405979|000|skin radiation necrosis
C1405979|000|lung radiation necrosis
C1405979|000|pulmonary radiation necrosis
C1405979|000|bone radiation necrosis
C1405979|000|mandibular radiation necrosis
C1405979|000|mandibular radionecrosis
C1405979|000|osteoradionecrosis
C1405979|000|radionecrosis of bone
C1405979|000|radionecrosis jaw
C1405979|000|radiation-induced bone necrosis
C1405979|000|soft tissue radionecrosis
C1405979|000|necrosis from rt
C1405979|000|necrosis from srs
C1405979|000|necrosis from radiosurgery
C1405979|000|necrosis from sbrt
C1405979|000|necrosis from gamma knife
C1405979|000|post-radiation necrotic change
C1405979|000|necrosis after irradiation
C1405979|000|necrosis following radiation therapy
C1405979|000|necrosis 2/2 radiation
C1405979|000|d/t rt necrosis
C1405979|000|post-xrt necrosis
C1405979|000|xrt necrosis
C1405979|000|ir necrosis
C1405979|000|necrosis s/p xrt
C1405979|000|necrosis d/t xrt
C1405979|000|necrosis post-xrt
C1405979|000|necrosis related to irradiation
C1405979|000|necrosis associated with radiation
C1405979|000|radiation damage with necrosis
C1405979|000|radiation-induced tissue necrosis
C1405979|000|tissue radionecrosis
C1405979|000|necrosis secondary to radiotherapy
C1405979|000|post-irradiation necrosis
C1405979|000|necrosis after beam therapy
C1405979|000|tissue death due to rt
C1405979|000|necrosis from therapeutic irradiation
C1405979|000|post-treatment necrosis (radiation)
C1405979|000|postradiosurgical necrosis
C1405979|000|sbrt-related necrosis
C1405979|000|srt-related necrosis
C1405979|000|stereotactic rt necrosis
C1405979|000|post-gamma knife necrosis
C1405979|000|gamma knife-induced necrosis
C1405979|000|irradiation effect necrosis
C1405979|000|irradiation-related necrosis
C1405979|000|necrosis subsequent to radiation
C1405979|000|necrosis subsequent to rt
C1405979|000|necrosis post radiotherapy
C1405979|000|necrosis after rt
C1405979|000|irradiation-associated necrosis
C1392786|000|cognitive dysfunction
C1392786|000|cognitive impairment
C1392786|000|cognitive decline
C1392786|000|cognitive deficits
C1392786|000|cognitive disturbance
C1392786|000|cognition impaired
C1392786|000|cognition changes
C1392786|000|altered cognition
C1392786|000|memory loss
C1392786|000|memory impairment
C1392786|000|forgetfulness
C1392786|000|short-term memory loss
C1392786|000|long-term memory loss
C1392786|000|confusion
C1392786|000|disorientation
C1392786|000|altered mental status
C1392786|000|ams
C1392786|000|encephalopathy
C1392786|000|delirium
C1392786|000|delirious
C1392786|000|acute mental status change
C1392786|000|fluctuating mental status
C1392786|000|clouded mentation
C1392786|000|mentation changes
C1392786|000|slowed mentation
C1392786|000|impaired executive function
C1392786|000|executive dysfunction
C1392786|000|difficulty concentrating
C1392786|000|concentration deficit
C1392786|000|decreased attention span
C1392786|000|attention deficit
C1392786|000|inattention
C1392786|000|impaired attention
C1392786|000|poor recall
C1392786|000|impaired recall
C1392786|000|impaired judgment
C1392786|000|judgment deficits
C1392786|000|difficulty making decisions
C1392786|000|reversible cognitive impairment
C1392786|000|irreversible cognitive impairment
C1392786|000|mild cognitive impairment
C1392786|000|mci
C1392786|000|dementia
C1392786|000|demented
C1392786|000|early-onset dementia
C1392786|000|late-onset dementia
C1392786|000|progressive cognitive decline
C1392786|000|vascular cognitive impairment
C1392786|000|vci
C1392786|000|ischemic cognitive impairment
C1392786|000|ischemic encephalopathy
C1392786|000|post-stroke cognitive changes
C1392786|000|stroke-related cognitive decline
C1392786|000|non-ischemic cognitive changes
C1392786|000|hypoxic encephalopathy
C1392786|000|hypoxic cognitive dysfunction
C1392786|000|chemo brain
C1392786|000|chemo-induced cognitive changes
C1392786|000|chemo-related cognitive impairment
C1392786|000|tumor-related cognitive change
C1392786|000|brain metastases cognitive effect
C1392786|000|radiation-induced cognitive decline
C1392786|000|amyloid-related cognitive impairment
C1392786|000|alzheimer's type changes
C1392786|000|ad-type dementia
C1392786|000|frontotemporal cognitive impairment
C1392786|000|ftd
C1392786|000|lewy body cognitive dysfunction
C1392786|000|dlb
C1392786|000|parkinson's-related cognitive change
C1392786|000|pd dementia
C1392786|000|ath-related cognitive dysfunction
C1392786|000|atherosclerotic cognitive impairment
C1392786|000|hypertensive encephalopathy
C1392786|000|hypertensive cognitive decline
C1392786|000|metabolic encephalopathy
C1392786|000|hepatic encephalopathy
C1392786|000|uremic encephalopathy
C1392786|000|sepsis-associated encephalopathy
C1392786|000|toxic-metabolic encephalopathy
C1392786|000|tme
C1392786|000|medication-related cognitive impairment
C1392786|000|polypharmacy-induced cognitive change
C1392786|000|sedative-induced confusion
C1392786|000|delirium due to meds
C1392786|000|alcohol-related cognitive dysfunction
C1392786|000|wernicke's encephalopathy
C1392786|000|korsakoff psychosis
C1392786|000|post-ictal confusion
C1392786|000|postictal cognitive changes
C1392786|000|epileptic cognitive dysfunction
C1392786|000|autoimmune encephalopathy
C1392786|000|paraneoplastic encephalopathy
C1392786|000|infectious encephalopathy
C1392786|000|hiv-associated neurocognitive disorder
C1392786|000|hand
C1392786|000|neurocognitive disorder
C1392786|000|ncd
C1392786|000|mild neurocognitive disorder
C1392786|000|major neurocognitive disorder
C1392786|000|cns dysfunction
C1392786|000|brain fog
C1392786|000|slowed cognition
C1392786|000|mental slowing
C1392786|000|mental clouding
C1392786|000|diminished cognition
C1392786|000|reduced cognitive capacity
C1392786|000|task management difficulty
C1392786|000|slowed thought process
C1392786|000|impaired thought process
C1392786|000|slowed reaction time
C1392786|000|reduced mental clarity
C1392786|000|mental dullness
C1392786|000|cognitive slowing
C1392786|000|depressive pseudodementia
C1392786|000|mood-related cognitive dysfunction
C1392786|000|psychosis-related cognitive change
C1392786|000|schizophrenia cognitive deficits
C1392786|000|bipolar cognitive dysfunction
C1392786|000|anoxic encephalopathy
C1392786|000|co poisoning cognitive effect
C1392786|000|encephalopathic
C1392786|000|icu psychosis
C1392786|000|hospital-acquired delirium
C1392786|000|postoperative cognitive dysfunction
C1392786|000|pocd
C1392786|000|sundowning
C1392786|000|pre-dementia state
C1392786|000|prodromal dementia
C1392786|000|subcortical dementia
C1392786|000|cortical dementia
C1392786|000|microvascular cognitive impairment
C1392786|000|subcortical ischemic cognitive change
C1392786|000|tbi cognitive deficits
C1392786|000|concussion cognitive changes
C1392786|000|blast injury cognitive change
C1392786|000|chronic traumatic encephalopathy
C1392786|000|cte
C1392786|000|huntington's cognitive impairment
C1392786|000|huntington's dementia
C1392786|000|wilson's disease cognitive change
C1392786|000|lyme neuroborreliosis cognitive effect
C1392786|000|post-covid cognitive dysfunction
C1392786|000|covid brain fog
C1392786|000|pasc cognitive change
C1392786|000|fatigue-related cognitive impairment
C1392786|000|sleep deprivation cognitive deficits
C1392786|000|obstructive sleep apnea cognitive change
C1392786|000|osa cognitive impairment
C1392786|000|drug-induced cognitive dysfunction
C1392786|000|thc-related cognitive change
C1392786|000|opioid-associated cognition change
C1392786|000|polytrauma cognitive deficits
C1392786|000|emotional distress-related cognition change
C1392786|000|adjustment disorder with cognitive symptoms
C1392786|000|adolescent cognitive changes
C1392786|000|geriatric cognitive decline
C1392786|000|aging-related cognitive change
C1392786|000|senile dementia
C1392786|000|senile cognitive changes
C1392786|000|mci-amnestic
C1392786|000|mci-nonamnestic
C1392786|000|attention/executive dysfunction
C1392786|000|language dysfunction
C1392786|000|praxis impairment
C1392786|000|visuospatial dysfunction
C1392786|000|agitation with cognitive impairment
C1392786|000|wandering with cognitive disorder
C1392786|000|anosognosia
C1392786|000|aphasia with cognitive decline
C1392786|000|agraphia/cognitive changes
C1392786|000|alexia/cognitive issues
C1392786|000|dysexecutive syndrome
C1392786|000|multifactorial cognitive impairment
C1392786|000|delirium superimposed on dementia
C0011206|000|delirium
C0011206|000|acute confusional state
C0011206|000|acs
C0011206|000|icu delirium
C0011206|000|hospital-acquired delirium
C0011206|000|acute brain failure
C0011206|000|subsyndromal delirium
C0011206|000|hyperactive delirium
C0011206|000|hypoactive delirium
C0011206|000|mixed delirium
C0011206|000|postoperative delirium
C0011206|000|post-op delirium
C0011206|000|post-anesthesia delirium
C0011206|000|emergence delirium
C0011206|000|agitated delirium
C0011206|000|toxic delirium
C0011206|000|metabolic delirium
C0011206|000|hepatic encephalopathy
C0011206|000|septic encephalopathy
C0011206|000|infectious delirium
C0011206|000|alcohol withdrawal delirium
C0011206|000|delirium tremens
C0011206|000|dts
C0011206|000|benzodiazepine withdrawal delirium
C0011206|000|drug-induced delirium
C0011206|000|chemo-induced delirium
C0011206|000|medication-induced delirium
C0011206|000|iatrogenic delirium
C0011206|000|icu psychosis
C0011206|000|sun-downing
C0011206|000|sundowning syndrome
C0011206|000|sundown syndrome
C0011206|000|acute encephalopathy
C0011206|000|fluctuating mental status
C0011206|000|waxing-waning mental status
C0011206|000|altered mental status
C0011206|000|ams
C0011206|000|mental status changes
C0011206|000|acute ams
C0011206|000|encephalopathic changes
C0011206|000|paranoid delirium
C0011206|000|delirious state
C0011206|000|clouded sensorium
C0011206|000|acute organic brain syndrome
C0011206|000|confusional syndrome
C0011206|000|toxic confusional state
C0011206|000|postictal confusion
C0011206|000|delirium superimposed on dementia
C0011206|000|delirium-on-dementia
C0011206|000|delirium of mixed etiology
C0011206|000|covid delirium
C0011206|000|hypoxemic delirium
C0011206|000|urosepsis delirium
C0011206|000|sepsis-associated delirium
C0011206|000|delirium due to uti
C0011206|000|delirium due to pneumonia
C0011206|000|perceptual disturbance
C0011206|000|psychomotor agitation
C0011206|000|psychomotor disturbance
C0011206|000|transient cognitive impairment
C0011206|000|transient delirium
C0011206|000|acute psychosis (delirium type)
C0011206|000|agitated confusion
C0011206|000|disorganized thinking
C0011206|000|attention deficit (acute)
C0011206|000|acute cognitive dysfunction
C0011206|000|perioperative delirium
C0011206|000|delirium of elderly
C0011206|000|delirium in dementia
C0011206|000|terminal delirium
C0011206|000|end-of-life delirium
C0011206|000|delirium in palliative care
C0011206|000|uremic encephalopathy
C0011206|000|hepatic delirium
C0011206|000|delirium secondary to infection
C0011206|000|delirium secondary to metabolic encephalopathy
C0011206|000|nonconvulsive status epilepticus with confusional state
C0011206|000|post-cardiac surgery delirium
C0011206|000|trauma-related delirium
C0011206|000|withdrawal delirium
C0011206|000|anticholinergic toxicity
C0011206|000|anticholinergic delirium
C0011206|000|delirium due to medication
C0011206|000|cns toxicity (delirium)
C0011206|000|delirium state
C0011206|000|delirium episode
C0011206|000|acute onset confusion
C0011206|000|delirious episode
C0011206|000|confusional episode
C0011206|000|acute cognitive change
C0011206|000|acute mental status change
C0011206|000|catatonic delirium
C0011206|000|poststroke delirium
C0011206|000|delirium due to stroke
C0011206|000|opiate-induced delirium
C0011206|000|pain control delirium
C0011206|000|cardiac surgery delirium
C0011206|000|anoxic delirium
C0011206|000|sleep deprivation delirium
C0011206|000|encephalopathic delirium
C0011206|000|toxic-metabolic encephalopathy
C0011206|000|endocrine delirium
C0011206|000|thyrotoxic encephalopathy
C0011206|000|thyroid storm delirium
C0011206|000|delirium due to cerebral hypoperfusion
C0011206|000|pediatric delirium
C0011206|000|delirium in children
C0011206|000|hepatic failure delirium
C0011206|000|delirium due to renal failure
C0011206|000|reversible encephalopathy
C0011206|000|wernicke's encephalopathy
C0011206|000|alcohol-related delirium
C0011206|000|stimulant-induced delirium
C0011206|000|delirium nos
C0011206|000|acute delirium episode
C0011206|000|delirium of advanced age
C0011206|000|delirium of critical illness
C0011206|000|delirium by dsm criteria
C0497327|000|dementia
C0497327|000|dem
C0497327|000|demented
C0497327|000|major neurocognitive disorder
C0497327|000|ncd
C0497327|000|chronic cognitive impairment
C0497327|000|cognitive decline
C0497327|000|cognitive dysfunction
C0497327|000|memory loss syndrome
C0497327|000|progressive cognitive decline
C0497327|000|senile dementia
C0497327|000|senile dem
C0497327|000|senile degeneration
C0497327|000|senile brain disease
C0497327|000|presenile dementia
C0497327|000|vascular dementia
C0497327|000|vad
C0497327|000|multi-infarct dementia
C0497327|000|arteriosclerotic dementia
C0497327|000|ischemic dementia
C0497327|000|post-stroke dementia
C0497327|000|alzheimer disease
C0497327|000|ad
C0497327|000|alzheimer's dementia
C0497327|000|alzheimer-type dementia
C0497327|000|mixed dementia
C0497327|000|dementia with lewy bodies
C0497327|000|dlb
C0497327|000|lewy body dementia
C0497327|000|frontotemporal dementia
C0497327|000|ftd
C0497327|000|pick disease
C0497327|000|pick's dementia
C0497327|000|subcortical dementia
C0497327|000|huntington dementia
C0497327|000|huntington's dementia
C0497327|000|hd dementia
C0497327|000|parkinsonian dementia
C0497327|000|parkinson's dementia
C0497327|000|pdd
C0497327|000|parkinsonism with dementia
C0497327|000|alcoholic dementia
C0497327|000|wernicke-korsakoff syndrome
C0497327|000|wks
C0497327|000|hiv-associated dementia
C0497327|000|had
C0497327|000|aids-dementia complex
C0497327|000|adc
C0497327|000|hiv dementia
C0497327|000|posttraumatic dementia
C0497327|000|traumatic dementia
C0497327|000|tbi-related dementia
C0497327|000|chronic traumatic encephalopathy
C0497327|000|cte
C0497327|000|creutzfeldt-jakob dementia
C0497327|000|creutzfeldt-jakob disease
C0497327|000|cjd
C0497327|000|prion dementia
C0497327|000|rapidly progressive dementia
C0497327|000|amyloid dementia
C0497327|000|autoimmune dementia
C0497327|000|hashimoto encephalopathy
C0497327|000|he dementia
C0497327|000|normal pressure hydrocephalus dementia
C0497327|000|nph dementia
C0497327|000|hydrocephalic dementia
C0497327|000|hepatic encephalopathy with dementia
C0497327|000|liver-related dementia
C0497327|000|hepatic dementia
C0497327|000|dialysis dementia
C0497327|000|uremic dementia
C0497327|000|metabolic dementia
C0497327|000|toxic dementia
C0497327|000|chemo-induced dementia
C0497327|000|chemotherapy-related cognitive impairment
C0497327|000|crci
C0497327|000|paraneoplastic dementia
C0497327|000|hypoxic-ischemic encephalopathy with dementia
C0497327|000|hie dementia
C0497327|000|hypoxic-ischemic dementia
C0497327|000|postanoxic dementia
C0497327|000|hypoglycemic dementia
C0497327|000|endocrine dementia
C0497327|000|thyroid dementia
C0497327|000|thyroid-related cognitive impairment
C0497327|000|syphilitic dementia
C0497327|000|neurosyphilis with dementia
C0497327|000|progressive paralytic dementia
C0497327|000|progressive general paralysis of the insane
C0497327|000|pgp
C0497327|000|dementia praecox
C0497327|000|madness
C0497327|000|organic brain syndrome
C0497327|000|obs
C0497327|000|chronic organic brain disorder
C0497327|000|cerebral degeneration
C0497327|000|brain failure
C0497327|000|global cognitive dysfunction
C0497327|000|general cognitive decline
C0497327|000|chronic encephalopathy
C0497327|000|irreversible cognitive decline
C0497327|000|idiopathic dementia
C0497327|000|primary dementia
C0497327|000|secondary dementia
C0497327|000|drug-induced cognitive impairment
C0497327|000|iatrogenic dementia
C0497327|000|nos dementia
C0497327|000|not otherwise specified dementia
C0497327|000|late-onset dementia
C0497327|000|early-onset dementia
C0497327|000|juvenile dementia
C0497327|000|mild dementia
C0497327|000|moderate dementia
C0497327|000|severe dementia
C0497327|000|advanced dementia
C0497327|000|terminal dementia
C0497327|000|rapid-onset dementia
C0497327|000|progressive dementia
C0497327|000|static dementia
C0497327|000|potentially reversible dementia
C0497327|000|irreversible dementia
C0497327|000|prodromal dementia
C0497327|000|amnestic syndrome
C0497327|000|amnestic disorder
C0497327|000|korsakoff dementia
C0497327|000|wernicke dementia
C0497327|000|non-ad dementia
C0497327|000|non-alzheimer dementia
C0497327|000|prion-related dementia
C0497327|000|motor neuron disease dementia
C0497327|000|als dementia
C0497327|000|amyotrophic lateral sclerosis dementia
C0497327|000|peripheral neuropathy with dementia
C0497327|000|diffuse lewy body disease
C0497327|000|familial dementia
C0497327|000|inherited dementia
C0497327|000|cerebral amyloid angiopathy-related dementia
C0497327|000|caa dementia
C0497327|000|cadasil-related dementia
C0497327|000|cadasil dementia
C0497327|000|notch3 dementia
C0497327|000|binswanger disease
C0497327|000|binswanger's dementia
C0497327|000|subcortical arteriosclerotic encephalopathy
C0497327|000|reversible dementia
C0497327|000|parkinson-plus dementia
C0497327|000|progressive supranuclear palsy dementia
C0497327|000|psp dementia
C0497327|000|corticobasal degeneration dementia
C0497327|000|cbd dementia
C0497327|000|dementia syndrome
C0497327|000|aphasic dementia
C0497327|000|semantic dementia
C0497327|000|logopenic dementia
C0497327|000|primary progressive aphasia
C0497327|000|ppa
C0497327|000|behavioral variant ftd
C0497327|000|bvftd
C0497327|000|semantic variant ppa
C0497327|000|nonfluent variant ppa
C0497327|000|nph cognitive impairment
C0497327|000|postinfectious dementia
C0497327|000|postmeningitic dementia
C0497327|000|herpes simplex encephalitis with dementia
C0497327|000|autoimmune encephalitis with dementia
C0497327|000|syndrome of dementia
C0497327|000|dementia-like syndrome
C0497327|000|mild cognitive impairment progressing to dementia
C0497327|000|mci progressing to dementia
C0497327|000|mci-to-dementia
C0497327|000|major ncd
C0497327|000|progressive memory loss
C0497327|000|intellectual deterioration
C0497327|000|generalized cognitive impairment
C0021125|000|impulsivity
C0021125|000|impulsive tendencies
C0021125|000|impulse control deficit
C0021125|000|impaired impulse control
C0021125|000|disinhibition
C0021125|000|disinhibited behavior
C0021125|000|behavioral disinhibition
C0021125|000|poor impulse control
C0021125|000|difficulty controlling impulses
C0021125|000|loss of impulse control
C0021125|000|acting on impulse
C0021125|000|compulsive urges
C0021125|000|compulsive actions
C0021125|000|lack of inhibition
C0021125|000|lack of self-control
C0021125|000|difficulty delaying gratification
C0021125|000|acts without thinking
C0021125|000|rash behavior
C0021125|000|impulsive acts
C0021125|000|impulsive responding
C0021125|000|impulsive actions
C0021125|000|impaired behavioral regulation
C0021125|000|reduced impulse control
C0021125|000|frontal lobe disinhibition
C0021125|000|frontal release
C0021125|000|auto-impulsive behavior
C0021125|000|impulsive decision-making
C0021125|000|poor behavioral inhibition
C0021125|000|diminished impulse control
C0021125|000|unrestrained behavior
C0021125|000|uncontrolled impulses
C0021125|000|lack of self-restraint
C0021125|000|executive dysfunction—impulsivity
C0021125|000|prefrontal syndrome—impulsivity
C0021125|000|hyperactivity—impulsivity
C0021125|000|bid (behavioral impulse dysregulation)
C0021125|000|icd (impulse control disorder)
C0021125|000|adhd-impulsivity
C0021125|000|addictive behavior
C0021125|000|mania—impulsivity
C0021125|000|manic impulsivity
C0021125|000|bpad—impulsivity
C0021125|000|tbi—disinhibition
C0021125|000|post-stroke impulsivity
C0021125|000|ischemic-frontal impulsivity
C0021125|000|nonischemic-frontal impulsivity
C0021125|000|frontotemporal disinhibition
C0021125|000|dementia-related impulsivity
C0021125|000|ad—disinhibition
C0021125|000|ftd—impulsive behavior
C0021125|000|vascular dementia—impulsive
C0021125|000|substance-induced disinhibition
C0021125|000|stimulant-induced impulsivity
C0021125|000|chemo-induced impulsivity
C0021125|000|iatrogenic impulsivity
C0021125|000|ssri-induced impulsivity
C0021125|000|ldopa-induced impulsivity
C0021125|000|pd—impulse control disorder
C0021125|000|pramipexole-induced impulsivity
C0021125|000|dopaminergic impulsivity
C0021125|000|ocd—impulsive symptoms
C0021125|000|borderline impulsivity
C0021125|000|antisocial behavior—impulsivity
C0021125|000|impulsive aggression
C0021125|000|impulsive self-harm
C0021125|000|parasuicidal impulsivity
C0021125|000|sib (self-injurious behavior)
C0021125|000|intermittent explosive episodes
C0021125|000|ied (intermittent explosive disorder)
C0021125|000|dysexecutive impulsivity
C0021125|000|executive function dysregulation
C0021125|000|cognitive impulsivity
C0021125|000|behavioral impulsivity
C0021125|000|motor impulsivity
C0021125|000|verbal impulsivity
C0021125|000|risk-taking behavior
C0021125|000|reckless behavior
C0021125|000|impulsive risk-taking
C0021125|000|failure to inhibit responses
C0021125|000|prepotent response disinhibition
C0021125|000|response inhibition deficit
C0021125|000|dysregulated behavior
C0021125|000|impulse-driven actions
C0021125|000|failure of behavioral restraint
C0021125|000|reward-driven impulsivity
C0021125|000|impulsive motor acts
C0021125|000|short latency responding
C0021125|000|failure to consider consequences
C0021125|000|acting without forethought
C0021125|000|split-second actions
C0021125|000|compromised self-regulation
C0021125|000|poor emotional regulation—impulsivity
C0021125|000|emotion-driven impulsivity
C0021125|000|ir (impulsive responding)
C0021125|000|irb (impulsive/reckless behavior)
C0021125|000|agitated impulsivity
C0021125|000|psychotic impulsivity
C0021125|000|bipolar impulsivity
C0021125|000|schizoaffective—impulsivity
C0021125|000|tic-related impulsivity
C0021125|000|impulsive outbursts
C0021125|000|impulsive speech
C0021125|000|loss of behavioral filter
C0021125|000|uninhibited actions
C0021125|000|loss of frontal lobe inhibition
C0021125|000|impulse dysregulation
C0021125|000|hyperimpulsivity
C0021125|000|pfc dysfunction—impulsivity
C0021125|000|corticobasal syndrome—impulsivity
C0021125|000|impulsive gambling
C0021125|000|compulsive spending—impulsivity
C0021125|000|hypersexuality—impulsivity
C0021125|000|substance binging—impulsivity
C0021125|000|poor delay of gratification
C0021125|000|impaired self-control
C0021125|000|urge-driven behavior
C0021125|000|ictal impulsivity
C0021125|000|seizure-related impulsivity
C0021125|000|irritable impulsivity
C0021125|000|impaired social inhibition
C0021125|000|reckless spending
C0021125|000|rage attacks
C0021125|000|sudden aggressive acts
C0021125|000|reckless driving
C0021125|000|impulsive shoplifting
C0021125|000|pathological impulsivity
C0021125|000|labile impulsivity
C0021125|000|transient disinhibition
C0021125|000|acute-onset disinhibition
C0021125|000|persistent impulsivity
C0021125|000|perseverative impulsivity
C0021125|000|interactive impulsivity
C0021125|000|adolescent impulsivity
C0021125|000|emotional disinhibition
C0021125|000|late-life impulsivity
C0021125|000|childhood impulsivity
C0021125|000|neurocognitive impulsivity
C0021125|000|neurobehavioral disinhibition
C0021125|000|postictal impulsivity
C0021125|000|parkinsonian impulsivity
C0021125|000|impulsive spending
C0021125|000|dysinhibition syndrome
C0021125|000|medication-induced impulsivity
C0021125|000|personality disorder—impulsivity
C0021125|000|impulsive suicidal behavior
C0021125|000|impulsive substance use
C0021125|000|alcohol-related impulsivity
C0021125|000|cns disorder—impulsivity
C0021125|000|chronic impulsivity
C0021125|000|executive system breakdown
C0021125|000|delay aversion
C0021125|000|frontal dysexecutive syndrome
C0021125|000|neurological impulsivity
C0021125|000|psychiatric impulsivity
C0021125|000|primary impulsivity
C0021125|000|secondary impulsivity
C0021125|000|disinhibition (psych/neuro)
C0021125|000|limbic impulsivity
C0021125|000|subcortical impulsivity
C0021125|000|posttraumatic impulsivity
C0021125|000|tbi—impulse control disorder
C0021125|000|impulsive sexual behavior
C0021125|000|shallow decision making
C0021125|000|prefrontal disinhibition
C0021125|000|hyperkinetic impulsivity
C0021125|000|impulsive binge eating
C0021125|000|psychostimulant-induced impulsivity
C0021125|000|parkinsonism—impulsivity
C0021125|000|ftd—behavioral disinhibition
C0021125|000|sud—impulsivity
C0021125|000|emotionally labile—impulsive
C0021125|000|mood-congruent impulsivity
C0021125|000|obsessive-impulsive behavior
C0021125|000|affective impulsivity
C0021125|000|paroxysmal impulsivity
C0021125|000|frontosubcortical impulsivity
C2748208|000|poor executive function
C2748208|000|impaired executive function
C2748208|000|executive dysfunction
C2748208|000|ef deficits
C2748208|000|executive impairment
C2748208|000|deficits in executive function
C2748208|000|executive fx deficits
C2748208|000|executive fx impairment
C2748208|000|dysfunctional executive function
C2748208|000|frontal lobe dysfunction
C2748208|000|frontal executive dysfunction
C2748208|000|executive cognitive deficit
C2748208|000|reduced executive capacity
C2748208|000|impaired ef
C2748208|000|ef impairment
C2748208|000|executive processing deficits
C2748208|000|decreased executive function
C2748208|000|frontal syndrome
C2748208|000|executive skill deficits
C2748208|000|executive control deficit
C2748208|000|impaired cognitive flexibility
C2748208|000|frontally-mediated impairment
C2748208|000|dysexecutive syndrome
C2748208|000|executive system dysfunction
C2748208|000|pfc impairment
C2748208|000|executive performance deficit
C2748208|000|executive control impairment
C2748208|000|cognitive control problems
C2748208|000|loss of executive function
C2748208|000|executive capacity loss
C2748208|000|impaired planning ability
C2748208|000|disorganized thinking
C2748208|000|working memory deficits
C2748208|000|frontal deficits
C2748208|000|frontostriatal dysfunction
C2748208|000|frontosubcortical impairment
C2748208|000|frontal-executive disorder
C2748208|000|frontal executive impairment
C2748208|000|executive fxn problems
C2748208|000|executive dysfunction d/t ad
C2748208|000|executive dysfunction in ftd
C2748208|000|vascular executive dysfunction
C2748208|000|executive dysfunction post-tbi
C2748208|000|executive dysfunction in schizophrenia
C2748208|000|executive dysfunction in mdd
C2748208|000|executive dysfunction in cte
C2748208|000|impaired executive network
C2748208|000|deficient executive processing
C2748208|000|decreased executive skills
C2748208|000|executive attention deficits
C2748208|000|frontal impairment
C2748208|000|executive d/o
C2748208|000|dysexecutive d/o
C2748208|000|frontal lobe syndrome
C2748208|000|impaired task switching
C2748208|000|dysregulated executive function
C2748208|000|impaired ability to plan
C2748208|000|organizing deficits
C2748208|000|sequencing deficits
C2748208|000|inhibition deficit
C2748208|000|problem-solving deficits
C2748208|000|impaired cognitive control
C2748208|000|executive problem
C2748208|000|executive planning difficulties
C2748208|000|loss of executive skills
C2748208|000|frontal circuit impairment
C2748208|000|executive fx difficulty
C2748208|000|executive fxn disruption
C2748208|000|impaired goal-directed behavior
C2748208|000|frontal-subcortical dysfunction
C2748208|000|frontally-based impairment
C2748208|000|pfc d/o
C2748208|000|executive domain impairment
C2748208|000|executive cognitive impairment
C2748208|000|impaired conceptualization
C2748208|000|executive network disruption
C2748208|000|executive impairment w/ vascular etiology
C2748208|000|executive syndrome
C2748208|000|executive control d/o
C2748208|000|abi-related executive dysfunction
C2748208|000|post-stroke executive deficits
C2748208|000|executive dysfunction in svd
C2748208|000|executive impairment secondary to frontal tumor
C2748208|000|executive fxn disorder
C2748208|000|executive processing impairment
C2748208|000|frontal executive deficits
C2748208|000|impaired set-shifting
C2748208|000|executive d/o nos
C2748208|000|executive fxn nos
C2748208|000|impairment in executive abilities
C2748208|000|executive pathway impairment
C2748208|000|dysexecutive pattern
C2748208|000|frontal dysexecutive syndrome
C2748208|000|frontal-executive deficits
C2748208|000|impaired response inhibition
C2748208|000|executive attention impairment
C2748208|000|pfc circuit dysfunction
C2748208|000|cognitive executive dysfunction
C2748208|000|defective executive function
C2748208|000|subcortical executive deficits
C2748208|000|frontal executive domain deficit
C2748208|000|disrupted executive function
C2748208|000|executive dysfunction s/p cva
C2748208|000|executive control failure
C2748208|000|executive dysfunction in adhd
C2748208|000|executive function weaknesses
C2748208|000|executive function disorder
C2748208|000|impaired higher-order control
C2748208|000|executive function abnormality
C2748208|000|executive function underfunction
C2748208|000|executive dysfunction nos
C2748208|000|frontal cognitive impairment
C2748208|000|dysexecutive impairment
C0751295|000|memory loss
C0751295|000|amnestic syndrome
C0751295|000|amnesia
C0751295|000|anterograde amnesia
C0751295|000|retrograde amnesia
C0751295|000|tga
C0751295|000|transient global amnesia
C0751295|000|short-term memory loss
C0751295|000|long-term memory loss
C0751295|000|memory impairment
C0751295|000|impaired memory
C0751295|000|cognitive impairment
C0751295|000|cognitive decline
C0751295|000|dementia
C0751295|000|ad
C0751295|000|alzheimer's disease
C0751295|000|vascular dementia
C0751295|000|multi-infarct dementia
C0751295|000|mild cognitive impairment
C0751295|000|mci
C0751295|000|age-associated memory impairment
C0751295|000|post-traumatic amnesia
C0751295|000|pta
C0751295|000|traumatic brain injury-related amnesia
C0751295|000|tbi-associated amnesia
C0751295|000|wernicke-korsakoff syndrome
C0751295|000|korsakoff amnesia
C0751295|000|alcohol-related amnesia
C0751295|000|chemo brain
C0751295|000|chemotherapy-induced cognitive impairment
C0751295|000|vascular amnestic syndrome
C0751295|000|hypoxic-ischemic memory loss
C0751295|000|stroke-related memory loss
C0751295|000|postictal amnesia
C0751295|000|epileptic amnesia
C0751295|000|tia-induced memory loss
C0751295|000|tia-related amnesia
C0751295|000|metabolic encephalopathy with memory loss
C0751295|000|encephalopathic memory disturbance
C0751295|000|delirium with impaired recall
C0751295|000|disorientation
C0751295|000|forgetfulness
C0751295|000|poor recall
C0751295|000|poor memory
C0751295|000|difficulty remembering
C0751295|000|loss of memory
C0751295|000|prion disease with memory loss
C0751295|000|creutzfeldt-jakob related memory loss
C0751295|000|frontotemporal dementia with memory deficits
C0751295|000|parkinson's dementia with memory impairment
C0751295|000|lewy body dementia with amnesia
C0751295|000|hiv-associated neurocognitive disorder with memory loss
C0751295|000|ancd
C0751295|000|ppa with memory involvement
C0751295|000|primary progressive aphasia with memory deficit
C0751295|000|mild amnestic changes
C0751295|000|remote memory loss
C0751295|000|recent memory loss
C0751295|000|febrile amnesia
C0751295|000|post-anoxic amnesia
C0751295|000|toxic encephalopathy with memory loss
C0751295|000|drug-induced amnesia
C0751295|000|medication-related memory loss
C0751295|000|anoxic brain injury-related memory loss
C0751295|000|limbic encephalitis with memory loss
C0751295|000|paraneoplastic limbic encephalitis with amnesia
C0751295|000|autoimmune encephalopathy with memory impairment
C0751295|000|hypoglycemic memory loss
C0751295|000|postictal confusion with amnesia
C0751295|000|infectious encephalopathy with amnesia
C0751295|000|hse memory loss
C0751295|000|herpes simplex encephalitis–related amnesia
C0751295|000|amnestic mild cognitive impairment
C0751295|000|amnestic mci
C0751295|000|global amnesia
C0751295|000|partial amnesia
C0751295|000|focal memory deficit
C0751295|000|subcortical amnesia
C0751295|000|hippocampal amnesia
C0751295|000|amygdalar memory loss
C0751295|000|psychiatric amnesia
C0751295|000|dissociative amnesia
C0751295|000|functional amnesia
C0751295|000|psychogenic amnesia
C0751295|000|hysterical amnesia
C0751295|000|trauma-induced memory loss
C0751295|000|concussion-related amnesia
C0751295|000|blackouts
C0751295|000|confabulatory memory disorder
C0751295|000|confabulation
C0751295|000|mild memory deficit
C0751295|000|significant memory impairment
C0751295|000|progressive memory loss
C0751295|000|chronic memory loss
C0751295|000|paroxysmal amnesia
C0751295|000|acute amnestic episode
C0751295|000|acute memory loss
C0751295|000|episodic memory loss
C0751295|000|semantic memory loss
C0751295|000|working memory deficit
C0751295|000|memory disturbance
C0751295|000|impaired recall
C0751295|000|impaired retention
C0751295|000|defective memory
C0751295|000|failing memory
C0751295|000|loss of retention
C0751295|000|historical amnesia
C0751295|000|anterograde deficit
C0751295|000|retrograde deficit
C0751295|000|ptsd-related amnesia
C0751295|000|stress-induced amnesia
C0751295|000|functional memory loss
C0751295|000|substance-induced memory loss
C0751295|000|prescribed medication-associated amnesia
C0751295|000|amnesia nos
C0751295|000|dementia-related memory loss
C0751295|000|cpm-related memory loss
C0751295|000|central pontine myelinolysis with amnesia
C0751295|000|tumor-related memory loss
C0751295|000|encephalopathic memory defect
C0751295|000|icu-acquired memory deficit
C0751295|000|icu delirium with impaired memory
C0751295|000|nonconvulsive status with amnesia
C0751295|000|nonconvulsive seizure with memory loss
C0751295|000|status epilepticus–related amnesia
C0751295|000|memory deficits
C0751295|000|recall difficulties
C0751295|000|early memory decline
C0751295|000|progressive amnestic disorder
C0751295|000|mild dementia with memory impairment
C0751295|000|mixed dementia with memory loss
C0751295|000|hypertensive encephalopathy with amnesia
C0751295|000|multi-etiology memory loss
C0751295|000|peripartum memory loss
C0751295|000|ppcm with memory impairment
C0751295|000|neurodegenerative memory loss
C0751295|000|amyloid-associated memory decline
C0751295|000|postinfectious memory loss
C0751295|000|hereditary amnesia
C0751295|000|genetic memory impairment
C0751295|000|autosomal dominant amnestic syndrome
C0751295|000|tauopathy with memory loss
C0751295|000|trauma-related memory impairment
C0751295|000|sedative-induced amnesia
C0751295|000|benzodiazepine-related amnesia
C0751295|000|anesthesia-associated amnesia
C0751295|000|anterograde memory deficit
C0751295|000|short-term amnesia
C0751295|000|long-term amnesia
C0751295|000|impaired long-term recall
C0751295|000|memory recall deficit
C0751295|000|subacute memory loss
C0751295|000|transient amnesia
C0751295|000|sudden-onset memory loss
C0751295|000|unexplained amnesia
C0751295|000|idiopathic memory loss
C0751295|000|unspecified amnesia
C0751295|000|attentional amnesia
C0751295|000|tia-induced amnesia
C0751295|000|silent infarct with memory loss
C0751295|000|nonischemic memory loss
C0751295|000|ischemic memory loss
C0751295|000|valvular memory loss
C0751295|000|hypertensive memory loss
C0751295|000|amyloid memory loss
C0751295|000|chemo-induced memory loss
C0751295|000|ppcm-associated memory loss
C0751295|000|tachycardia-induced memory loss
C0751295|000|myocarditis-associated memory loss
C0233794|000|memory impairment
C0233794|000|memory loss
C0233794|000|impaired memory
C0233794|000|amnestic syndrome
C0233794|000|amnesia
C0233794|000|memory dysfunction
C0233794|000|decreased memory
C0233794|000|poor memory
C0233794|000|short-term memory loss
C0233794|000|long-term memory loss
C0233794|000|stm loss
C0233794|000|ltm loss
C0233794|000|anterograde amnesia
C0233794|000|retrograde amnesia
C0233794|000|transient global amnesia
C0233794|000|tga
C0233794|000|transient amnesia
C0233794|000|memory deficit
C0233794|000|cognitive impairment
C0233794|000|ci
C0233794|000|memory disturbance
C0233794|000|deficit of recall
C0233794|000|recall impairment
C0233794|000|encoding deficit
C0233794|000|retrieval deficit
C0233794|000|executive memory dysfunction
C0233794|000|working memory impairment
C0233794|000|working memory deficit
C0233794|000|wmi
C0233794|000|impaired recall
C0233794|000|impaired retention
C0233794|000|dementia
C0233794|000|early dementia
C0233794|000|amnestic mci
C0233794|000|amci
C0233794|000|mci
C0233794|000|mild cognitive impairment
C0233794|000|vuci (vascular unrelated cognitive impairment)
C0233794|000|vci (vascular cognitive impairment)
C0233794|000|post-stroke memory loss
C0233794|000|ischemic memory loss
C0233794|000|vascular memory deficit
C0233794|000|nonischemic memory loss
C0233794|000|hypoxic memory impairment
C0233794|000|hypoxic brain injury with memory loss
C0233794|000|postencephalitic memory loss
C0233794|000|encephalopathic memory deficit
C0233794|000|tbi memory loss
C0233794|000|post-concussive amnesia
C0233794|000|concussion-related memory loss
C0233794|000|chemotherapy-induced memory impairment
C0233794|000|chemo brain
C0233794|000|radiation-induced memory deficit
C0233794|000|alcohol-related memory impairment
C0233794|000|wernicke-korsakoff amnesia
C0233794|000|wks
C0233794|000|thiamine deficiency–related memory loss
C0233794|000|alzheimer's-related memory loss
C0233794|000|ad-associated memory loss
C0233794|000|ftd memory loss
C0233794|000|frontotemporal dementia memory deficit
C0233794|000|pca memory impairment
C0233794|000|posterior cortical atrophy with memory loss
C0233794|000|lewy body dementia–associated memory loss
C0233794|000|lbd memory loss
C0233794|000|parkinson's with memory impairment
C0233794|000|pd memory deficit
C0233794|000|multiple sclerosis with memory loss
C0233794|000|ms-related memory impairment
C0233794|000|huntington’s chorea with memory loss
C0233794|000|amyloid-related memory impairment
C0233794|000|neurodegenerative memory loss
C0233794|000|iatrogenic memory deficit
C0233794|000|medication-related memory loss
C0233794|000|benzo-induced memory loss
C0233794|000|steroid-induced cognitive impairment
C0233794|000|psychiatric memory loss
C0233794|000|ptsd-related memory gap
C0233794|000|depressive pseudodementia
C0233794|000|anxiety-related memory impairment
C0233794|000|stress-induced memory deficit
C0233794|000|age-associated memory impairment
C0233794|000|aami
C0233794|000|presbycognitive change
C0233794|000|elderly memory decline
C0233794|000|mild memory decline
C0233794|000|subjective memory complaint
C0233794|000|forgetfulness
C0233794|000|recent memory deficit
C0233794|000|remote memory deficit
C0233794|000|remote memory impairment
C0233794|000|recognition impairment
C0233794|000|impaired knowledge retention
C0233794|000|deficient recall
C0233794|000|blackout (memory)
C0233794|000|global amnesia
C0233794|000|functional amnesia
C0233794|000|psychogenic amnesia
C0233794|000|dissociative amnesia
C0233794|000|hysterical amnesia
C0233794|000|traumatic amnesia
C0233794|000|reversible memory impairment
C0233794|000|irreversible memory impairment
C0233794|000|progressive memory loss
C0233794|000|episodic memory loss
C0233794|000|semantic memory loss
C0233794|000|immediate memory deficit
C0233794|000|delayed recall loss
C0233794|000|impaired new learning
C0233794|000|learning disability (acquired)
C0233794|000|impaired memory acquisition
C0233794|000|anterograde deficit
C0233794|000|retrograde deficit
C0233794|000|amnesic syndrome
C0233794|000|drug-induced amnesia
C0233794|000|toxic encephalopathy with memory loss
C0233794|000|metabolic encephalopathy with memory impairment
C0233794|000|autoimmune encephalitis–associated memory loss
C0233794|000|limbic encephalitis–associated memory loss
C0233794|000|temporal lobe memory deficit
C0233794|000|frontal lobe memory deficit
C0233794|000|medial temporal amnesia
C0233794|000|devastating memory loss
C0233794|000|attentional memory deficit
C0233794|000|ppcm-related cognitive deficit
C0233794|000|post-infectious cognitive impairment
C0233794|000|covid-related cognitive impairment
C0233794|000|long covid memory issues
C0233794|000|hiv-associated neurocognitive memory loss
C0233794|000|hand
C0233794|000|cjd memory loss
C0233794|000|prion-related memory deficit
C0233794|000|chronic memory loss
C0233794|000|acute memory loss
C0233794|000|subacute memory loss
C0233794|000|abrupt memory deficit
C0233794|000|persistent memory impairment
C0233794|000|fluctuating memory impairment
C0233794|000|paraneoplastic-related memory deficit
C0233794|000|seizure-associated amnesia
C0233794|000|postictal amnesia
C0233794|000|postictal confusion with memory loss
C0233794|000|epileptic amnesia
C0233794|000|epilepsy-related memory impairment
C0233794|000|temporal lobe epilepsy amnesia
C0233794|000|tle-associated memory loss
C0233794|000|atrial fibrillation–related memory loss
C0233794|000|af-related cognitive deficit
C0233794|000|hypertensive memory deficit
C0233794|000|cardiac memory loss
C0233794|000|chf-related memory impairment
C0233794|000|heart failure–associated cognitive impairment
C0233794|000|tachycardia-induced cognitive dysfunction
C0233794|000|tci-related memory loss
C0233794|000|neuropathic memory deficit
C0233794|000|cortical memory impairment
C0233794|000|subcortical memory impairment
C0233794|000|hie-related memory loss
C0233794|000|hypoxic-ischemic encephalopathy with memory loss
C0233794|000|hypoperfusion-related cognitive deficit
C0233794|000|dialysis dementia
C0233794|000|renal failure-related memory loss
C0233794|000|hepatic encephalopathy with memory deficit
C0233794|000|liver failure–related cognitive disorder
C0233794|000|systemic illness–related memory impairment
C0233794|000|delirium-associated amnesia
C0233794|000|icu-related memory deficit
C0233794|000|post-surgical memory loss
C0233794|000|perioperative amnesia
C0233794|000|critical illness–associated cognitive impairment
C0233407|000|disoriented
C0233407|000|disorientation
C0233407|000|ams
C0233407|000|altered mental status
C0233407|000|confusion
C0233407|000|confused
C0233407|000|delirium
C0233407|000|delirious
C0233407|000|mental status changes
C0233407|000|acute confusional state
C0233407|000|waxing and waning mental status
C0233407|000|disorganized thought process
C0233407|000|disorganized thought
C0233407|000|incoherent
C0233407|000|encephalopathy
C0233407|000|acute encephalopathy
C0233407|000|lethargy
C0233407|000|obtunded
C0233407|000|clouded sensorium
C0233407|000|mental clouding
C0233407|000|senile confusion
C0233407|000|acute mental status change
C0233407|000|altered level of consciousness
C0233407|000|near-syncope with confusion
C0233407|000|post-ictal confusion
C0233407|000|toxic-metabolic encephalopathy
C0233407|000|confusional state
C0233407|000|transient confusion
C0233407|000|acute organic brain syndrome
C0233407|000|disorientation to time
C0233407|000|disorientation to place
C0233407|000|disorientation to person
C0233407|000|chrono-disorientation
C0233407|000|spatial disorientation
C0233407|000|person-place-time disorientation
C0233407|000|aox1
C0233407|000|aox2
C0233407|000|aox3
C0233407|000|not aox3
C0233407|000|not alert and oriented
C0233407|000|poor orientation
C0233407|000|oriented x1
C0233407|000|oriented x2
C0233407|000|oriented x0
C0233407|000|diminished awareness
C0233407|000|no orientation
C0233407|000|stuporous
C0233407|000|disoriented behavior
C0233407|000|mental fog
C0233407|000|altered sensorium
C0233407|000|disoriented to surroundings
C0233407|000|cognitive dysfunction
C0233407|000|cognitive impairment
C0233407|000|acute mental confusion
C0233407|000|waxing/waning orientation
C0233407|000|episodes of confusion
C0233407|000|vague mentation
C0233407|000|inattentive
C0233407|000|memory lapse with confusion
C0233407|000|icu delirium
C0233407|000|hosp. delirium
C0233407|000|sun-downing
C0233407|000|sundowning
C0233407|000|critical illness encephalopathy
C0233407|000|hepatic encephalopathy
C0233407|000|uremic encephalopathy
C0233407|000|metabolic encephalopathy
C0233407|000|hypoxic encephalopathy
C0233407|000|septic encephalopathy
C0233407|000|postictal state
C0233407|000|confusional episode
C0233407|000|transient disorientation
C0233407|000|altered awareness
C0233407|000|impaired orientation
C0233407|000|o/e: disoriented
C0233407|000|aox1 (person)
C0233407|000|aox1 (place)
C0233407|000|aox1 (time)
C0233407|000|unoriented
C0233407|000|not oriented
C0233407|000|losing orientation
C0233407|000|fluctuating mental status
C0233407|000|acute onset confusion
C0233407|000|dementia-related confusion
C0233407|000|psychotic disorganization
C0233407|000|mental status waxing/waning
C0233407|000|short-term confusion
C0233407|000|periodic confusion
C0233407|000|post-operative confusion
C0233407|000|icu psychosis
C0233407|000|post-op delirium
C0233407|000|chemotherapy-induced delirium
C0233407|000|drug-induced confusion
C0233407|000|intoxication delirium
C0233407|000|withdrawal-related confusion
C0233407|000|alcoholic encephalopathy
C0233407|000|wernicke's encephalopathy
C0233407|000|delirium tremens
C0233407|000|tachycardia-induced confusion
C0233407|000|sepsis-induced ams
C0233407|000|infection-related altered mentation
C0233407|000|ppcm-related ams
C0233407|000|myocarditis delirium
C0233407|000|ischemic encephalopathy
C0233407|000|stroke-related confusion
C0233407|000|tia-related ams
C0233407|000|vascular dementia w/ confusion
C0233407|000|valvular disease ams
C0233407|000|hypertensive encephalopathy
C0233407|000|amyloid encephalopathy
C0233407|000|hypoglycemia with confusion
C0233407|000|hyperglycemic confusion
C0233407|000|dka-related ams
C0233407|000|hhs with disorientation
C0233407|000|hypercapnic encephalopathy
C0233407|000|co2 narcosis
C0233407|000|hypoxemic confusion
C0233407|000|anoxic encephalopathy
C0233407|000|thiamine-deficiency encephalopathy
C0233407|000|nonconvulsive status ams
C0233407|000|paraneoplastic encephalopathy
C0233407|000|tumor-related confusion
C0233407|000|brain metastasis ams
C0233407|000|space-occupying lesion ams
C0233407|000|subdural hematoma with confusion
C0233407|000|sah with disorientation
C0233407|000|traumatic brain injury ams
C0233407|000|mild cognitive impairment with confusion
C0233407|000|multifactorial ams
C0233407|000|confusional syndrome
C0233407|000|encephalopathic state
C0233407|000|organic brain syndrome
C0233407|000|momentary confusion
C0233407|000|low arousal state
C0233407|000|poor mentation
C0233407|000|encephalopathic changes
C0233407|000|delayed mentation
C0233407|000|nonresponsive with confusion
C0233407|000|unresponsive with confusion
C0233407|000|somnolent
C0233407|000|stupor with disorientation
C0233407|000|not alert
C0233407|000|disorganized mentation
C0233407|000|psychomotor disorientation
C0233407|000|cerebral dysfunction
C0233407|000|disoriented to environment
C0233407|000|no orientation to date
C0233407|000|no orientation to location
C0233407|000|acute confusion state
C0233407|000|hyperactive delirium
C0233407|000|hypoactive delirium
C0233407|000|mixed delirium
C0233407|000|fluctuating orientation
C0233407|000|confused on exam
C0233407|000|disoriented on assessment
C0233407|000|not oriented on exam
C0233407|000|o/e: confused
C0233407|000|patient confused
C0233407|000|pt confused
C0233407|000|pt disoriented
C0233407|000|aox0
C0233407|000|unaware of time/place
C0233407|000|disorientation to situation
C0233407|000|not oriented to time
C0233407|000|not oriented to place
C0233407|000|not oriented to self
C0233407|000|not oriented to situation
C0233407|000|orientation deficit
C0233407|000|aox
C0233407|000|impaired consciousness
C0233407|000|poor cognition
C0233407|000|acute altered consciousness
C0233407|000|mental slowing
C0233407|000|ams of unclear etiology
C0233407|000|global confusion
C0233407|000|cerebral confusion
C0233407|000|organic confusion
C0233407|000|cns dysfunction with confusion
C0233407|000|mental status alteration
C0233407|000|loss of orientation
C0233407|000|labile orientation
C0233407|000|impaired mentation
C0233407|000|not ao
C0233407|000|disturbed consciousness
C0015676|000|mental fatigue
C0015676|000|cognitive fatigue
C0015676|000|cognitive exhaustion
C0015676|000|cognitive weariness
C0015676|000|psychic fatigue
C0015676|000|psychic exhaustion
C0015676|000|psychic weariness
C0015676|000|neurofatigue
C0015676|000|neurocognitive fatigue
C0015676|000|mental exhaustion
C0015676|000|mental weariness
C0015676|000|mental tiredness
C0015676|000|cognitive tiredness
C0015676|000|psychological fatigue
C0015676|000|brain fatigue
C0015676|000|brain fog
C0015676|000|brain tiredness
C0015676|000|mental sluggishness
C0015676|000|decreased mental stamina
C0015676|000|neural fatigue
C0015676|000|cognitive slowing
C0015676|000|decreased cognitive endurance
C0015676|000|decreased concentration endurance
C0015676|000|loss of mental stamina
C0015676|000|reduced cognitive capacity
C0015676|000|subjective cognitive fatigue
C0015676|000|cerebral fatigue
C0015676|000|cortical fatigue
C0015676|000|chemo brain
C0015676|000|chemo-induced cognitive fatigue
C0015676|000|chemo-related brain fog
C0015676|000|crf (cancer-related fatigue)
C0015676|000|crcf (cancer-related cognitive fatigue)
C0015676|000|ms-related cognitive fatigue
C0015676|000|stroke-related mental fatigue
C0015676|000|ischemic cognitive fatigue
C0015676|000|nonischemic mental fatigue
C0015676|000|tbi-related mental fatigue
C0015676|000|postconcussive fatigue
C0015676|000|neurological fatigue
C0015676|000|als-related cognitive fatigue
C0015676|000|pd-related cognitive fatigue
C0015676|000|dementia-related fatigue
C0015676|000|depression-related fatigue
C0015676|000|post-stroke cognitive fatigue
C0015676|000|cfs-related mental fatigue
C0015676|000|chronic fatigue syndrome mental exhaustion
C0015676|000|primary fatigue of ms
C0015676|000|encephalopathic fatigue
C0015676|000|paraneoplastic fatigue
C0015676|000|autoimmune encephalitis cognitive fatigue
C0015676|000|ra-related mental fatigue
C0015676|000|lupus-related cognitive fatigue
C0015676|000|post-viral fatigue
C0015676|000|long covid brain fog
C0015676|000|pasc cognitive fatigue
C0015676|000|mental lassitude
C0015676|000|mental depletion
C0015676|000|attention fatigue
C0015676|000|executive fatigue
C0015676|000|decision fatigue
C0015676|000|sustained attention impairment
C0015676|000|mental stamina loss
C0015676|000|cognitive burnout
C0015676|000|mental burnout
C0015676|000|neuropsychiatric fatigue
C0015676|000|postictal fatigue
C0015676|000|post-seizure cognitive fatigue
C0015676|000|fibro fog
C0015676|000|fibromyalgia-related cognitive fatigue
C0015676|000|psychiatric fatigue
C0015676|000|schizophrenia-related cognitive fatigue
C0015676|000|bipolar-related cognitive fatigue
C0015676|000|ptsd-related cognitive fatigue
C0015676|000|csf (chronic symptom fatigue)
C0015676|000|chronic illness fatigue
C0015676|000|pots-related cognitive fatigue
C0015676|000|orthostatic cognitive fatigue
C0015676|000|dysautonomia fatigue
C0015676|000|anemia-related mental fatigue
C0015676|000|metabolic fatigue
C0015676|000|liver disease-related mental fatigue
C0015676|000|ckd-related cognitive fatigue
C0015676|000|dialysis-related cognitive fatigue
C0015676|000|hypothyroidism-related cognitive fatigue
C0015676|000|sle mental fatigue
C0015676|000|immune-mediated cognitive fatigue
C0015676|000|cancer brain fog
C0015676|000|brain fatigue syndrome
C0015676|000|postviral fatigue syndrome
C0015676|000|vaccination-related cognitive fatigue
C0015676|000|viral encephalitis-related fatigue
C0015676|000|substance-induced mental fatigue
C0015676|000|medication-induced cognitive fatigue
C0015676|000|drug-induced cognitive fatigue
C0015676|000|cognitive malaise
C0015676|000|nonrestorative cognitive fatigue
C0015676|000|fatigued cognition
C0015676|000|overtired mental state
C0015676|000|prolonged cognitive fatigue
C0015676|000|prolonged mental exhaustion
C0015676|000|work-related mental fatigue
C0015676|000|post-work mental exhaustion
C0015676|000|shift work-related mental fatigue
C0015676|000|vhf (viral hemorrhagic fever) related fatigue
C0015676|000|covid-19 related brain fog
C0015676|000|fatigue of central origin
C0015676|000|central fatigue
C0015676|000|pervasive cognitive fatigue
C0015676|000|psychomotor slowing
C0015676|000|cognitive inefficiency
C0015676|000|mental inefficiency
C0015676|000|cognitive drain
C0015676|000|mental drain
C0015676|000|cognitive depletion
C0015676|000|ptf (post-traumatic fatigue)
C0015676|000|fatigue nos
C0015676|000|subjective mental fatigue
C0015676|000|subjective brain fog
C0015676|000|reduced cognitive throughput
C0015676|000|cognitive wearout
C0015676|000|cognitive clouding
C0015676|000|mental fog
C0015676|000|decreased processing speed
C0015676|000|information processing fatigue
C0015676|000|executive function fatigue
C0015676|000|mental lethargy
C0015676|000|cognitive lethargy
C0015676|000|mental clouding
C0015676|000|cognitive cloudiness
C0015676|000|brain exhaustion
C0015676|000|mental enervation
C0015676|000|cognitive enervation
C0015676|000|loss of mental acuity
C0015676|000|decreased alertness
C0015676|000|sustained attention fatigue
C0015676|000|prolonged attentional fatigue
C0015676|000|prolonged vigilance fatigue
C0015676|000|vigilance decrement
C0015676|000|alertness decline
C0015676|000|delayed mental response
C0015676|000|mental processing delay
C0015676|000|cortical exhaustion
C0015676|000|frontal fatigue
C0015676|000|frontosubcortical fatigue
C0015676|000|psychogenic fatigue
C0015676|000|psychological exhaustion
C0015676|000|psychological tiredness
C0015676|000|occupational cognitive fatigue
C0015676|000|occupational brain fatigue
C0015676|000|task-related mental fatigue
C0015676|000|task-induced fatigue
C0015676|000|workload-related cognitive fatigue
C0015676|000|shiftwork fatigue
C0015676|000|driver fatigue (mental)
C0015676|000|operator mental fatigue
C0015676|000|performance fatigue
C0015676|000|mental overexertion
C0015676|000|cerebral exhaustion
C0015676|000|cognitive slowing syndrome
C0015676|000|effort fatigue
C0015676|000|expended cognitive reserves
C0015676|000|decreased cognitive reserves
C0015676|000|mental performance decrement
C0015676|000|mental function decrement
C0015676|000|ppcs-related fatigue
C0015676|000|post-tia cognitive fatigue
C0015676|000|hiv-associated neurocognitive fatigue
C0015676|000|aids-related cognitive fatigue
C0015676|000|immunotherapy-related brain fog
C0015676|000|antiviral-induced cognitive fatigue
C0015676|000|anticholinergic-related cognitive fatigue
C0015676|000|steroid-related cognitive fatigue
C0015676|000|anti-epileptic-induced cognitive fatigue
C0015676|000|antipsychotic-related cognitive fatigue
C0015676|000|depressogenic fatigue
C0015676|000|icu-related cognitive fatigue
C0015676|000|post-icu fatigue
C0015676|000|post-hospitalization mental fatigue
C0015676|000|sleep deprivation-related mental fatigue
C0015676|000|insomnia-related cognitive fatigue
C0015676|000|sleep disorder mental fatigue
C0015676|000|hypersomnia mental fatigue
C0015676|000|shiftwork disorder-related mental fatigue
C0015676|000|disrupted circadian cognitive fatigue
C0015676|000|nocturnal cognitive fatigue
C0015676|000|daytime cognitive fatigue
C0029227|000|delirium
C0029227|000|acute confusional state
C0029227|000|acute brain syndrome
C0029227|000|acute encephalopathy
C0029227|000|icu psychosis
C0029227|000|toxic encephalopathy
C0029227|000|substance-induced delirium
C0029227|000|alcohol withdrawal delirium
C0029227|000|dts
C0029227|000|delirium tremens
C0029227|000|hyperactive delirium
C0029227|000|hypoactive delirium
C0029227|000|mixed delirium
C0029227|000|dementia
C0029227|000|major neurocognitive disorder
C0029227|000|minor neurocognitive disorder
C0029227|000|neurocognitive disorder nos
C0029227|000|ncd
C0029227|000|primary degenerative dementia
C0029227|000|senile dementia
C0029227|000|presenile dementia
C0029227|000|senile cortical degeneration
C0029227|000|multi-infarct dementia
C0029227|000|mid
C0029227|000|vascular dementia
C0029227|000|vad
C0029227|000|ischemic vascular dementia
C0029227|000|nonischemic dementia
C0029227|000|subcortical dementia
C0029227|000|frontotemporal dementia
C0029227|000|ftd
C0029227|000|pick's disease
C0029227|000|lewy body dementia
C0029227|000|lbd
C0029227|000|parkinson’s disease dementia
C0029227|000|pdd
C0029227|000|alzheimer’s disease
C0029227|000|ad
C0029227|000|alzheimers type dementia
C0029227|000|dementia with behavioral disturbance
C0029227|000|dementia with psychosis
C0029227|000|dementia with delusions
C0029227|000|dementia with agitation
C0029227|000|dementia with depression
C0029227|000|aids dementia complex
C0029227|000|hiv-associated dementia
C0029227|000|hivd
C0029227|000|chemo-induced cognitive impairment
C0029227|000|chemotherapy-related cognitive dysfunction
C0029227|000|chemo brain
C0029227|000|alcohol-related dementia
C0029227|000|wernicke-korsakoff syndrome
C0029227|000|wks
C0029227|000|korsakoff dementia
C0029227|000|wernicke’s encephalopathy
C0029227|000|normal pressure hydrocephalus
C0029227|000|nph
C0029227|000|post-stroke dementia
C0029227|000|postinfectious dementia
C0029227|000|pandas encephalopathy
C0029227|000|creutzfeldt-jakob disease
C0029227|000|prion disease dementia
C0029227|000|huntington’s disease dementia
C0029227|000|hd dementia
C0029227|000|rapidly progressive dementia
C0029227|000|progressive supranuclear palsy dementia
C0029227|000|depression-related cognitive impairment
C0029227|000|pseudo-dementia
C0029227|000|amnestic disorder
C0029227|000|amnestic syndrome
C0029227|000|amnestic mci
C0029227|000|anoxic brain injury dementia
C0029227|000|hypoxic-ischemic encephalopathy
C0029227|000|down syndrome dementia
C0029227|000|ds dementia
C0029227|000|mild cognitive impairment
C0029227|000|mci
C0029227|000|age-related cognitive decline
C0029227|000|cognitive disorder nos
C0029227|000|organic brain syndrome
C0029227|000|obs
C0029227|000|organic mental disorder
C0029227|000|omd
C0029227|000|cognitive dysfunction
C0029227|000|cognitive decline
C0029227|000|chronic confusional state
C0029227|000|global cognitive impairment
C0029227|000|memory loss
C0029227|000|short-term memory loss
C0029227|000|long-term memory loss
C0029227|000|executive dysfunction
C0029227|000|aphasic dementia
C0029227|000|primary progressive aphasia
C0029227|000|semantic dementia
C0029227|000|logopenic progressive aphasia
C0029227|000|agrammatic aphasia
C0029227|000|cadasil dementia
C0029227|000|amyloid angiopathy-related dementia
C0029227|000|posterior cortical atrophy
C0029227|000|binswanger's disease
C0029227|000|thalamic dementia
C0029227|000|corticobasal degeneration dementia
C0029227|000|cbd dementia
C0029227|000|marchiafava-bignami disease
C0029227|000|menstrual-related cognitive changes
C0029227|000|steroid-induced cognitive dysfunction
C0029227|000|medication-induced encephalopathy
C0029227|000|paraneoplastic encephalopathy
C0029227|000|autoimmune encephalopathy
C0029227|000|anti-nmda receptor encephalitis
C0029227|000|syphilitic dementia
C0029227|000|neurosyphilis dementia
C0029227|000|wilson’s disease dementia
C0029227|000|copper-related cognitive disorder
C0029227|000|b12 deficiency dementia
C0029227|000|hypothyroid dementia
C0029227|000|hypoglycemic encephalopathy
C0029227|000|hypoparathyroidism cognitive dysfunction
C0029227|000|hypercalcemia cognitive impairment
C0029227|000|postictal confusion
C0029227|000|chronic traumatic encephalopathy
C0029227|000|cte
C0029227|000|ptsd-related cognitive disorder
C0029227|000|cognitive impairment nos
C0029227|000|transient global amnesia
C0029227|000|tga
C0029227|000|fahr's syndrome dementia
C0029227|000|basal ganglia dementia
C0029227|000|epileptic encephalopathy
C0029227|000|retrospective amnesia
C0029227|000|anterograde amnesia
C0029227|000|retrograde amnesia
C0029227|000|secondary dementia
C0029227|000|delirious mania
C0029227|000|steroid psychosis
C0029227|000|icu delirium
C0029227|000|withdrawal delirium
C0029227|000|metabolic encephalopathy
C0029227|000|hepatic encephalopathy
C0029227|000|uremic encephalopathy
C0029227|000|dialysis dementia
C0029227|000|dialysis encephalopathy
C0029227|000|hypoxic encephalopathy
C0029227|000|hypoxic-ischemic brain injury
C0029227|000|acute memory loss
C0029227|000|psychosis with cognitive decline
C0029227|000|behavioral variant dementia
C0029227|000|semantic variant primary progressive aphasia
C0029227|000|nonfluent variant primary progressive aphasia
C0029227|000|progressive nonfluent aphasia
C0029227|000|alzheimer-type psychosis
C0029227|000|mild ncd
C0029227|000|major ncd
C0029227|000|cognitive disorder due to trauma
C0029227|000|postconcussive syndrome cognitive deficit
C0029227|000|residual cognitive deficits
C0029227|000|ppcm cognitive disorder
C0029227|000|postpartum cognitive impairment
C0029227|000|peripartum cognitive disorder
C0029227|000|tachycardia-induced encephalopathy
C0029227|000|valvular-related dementia
C0029227|000|amyloid-related cognitive impairment
C0029227|000|toxic-metabolic encephalopathy
C0029227|000|dementia nos
C0029227|000|senile ncd
C0029227|000|mixed ncd
C0029227|000|age-associated memory impairment
C0029227|000|aami
C0029227|000|cortical dementia
C0029227|000|subcortical cognitive disorder
C0029227|000|ischemic encephalopathy
C0029227|000|hypertensive encephalopathy
C0029227|000|cadasil cognitive impairment
C0029227|000|binswanger type ncd
C0029227|000|cerebral amyloid angiopathy cognitive dysfunction
C0009676|000|confusion
C0009676|000|confused
C0009676|000|ams
C0009676|000|altered mental status
C0009676|000|acute confusion
C0009676|000|delirium
C0009676|000|encephalopathy
C0009676|000|acute encephalopathy
C0009676|000|subacute confusion
C0009676|000|disoriented
C0009676|000|disorientation
C0009676|000|impaired consciousness
C0009676|000|clouded sensorium
C0009676|000|impaired awareness
C0009676|000|decreased alertness
C0009676|000|impaired mentation
C0009676|000|drowsy
C0009676|000|obtunded
C0009676|000|lethargic
C0009676|000|waxing/waning level of consciousness
C0009676|000|inattentive
C0009676|000|difficulty following commands
C0009676|000|mental status change
C0009676|000|acute mental status change
C0009676|000|cognitive dysfunction
C0009676|000|cognitive disturbance
C0009676|000|delirious
C0009676|000|somnolent
C0009676|000|fluctuating mental status
C0009676|000|with confusion
C0009676|000|episodes of confusion
C0009676|000|disorganized thinking
C0009676|000|impaired thought process
C0009676|000|slowed thought process
C0009676|000|slowed cognition
C0009676|000|stuporous
C0009676|000|coma
C0009676|000|minimally responsive
C0009676|000|encephalopathic
C0009676|000|toxic/metabolic encephalopathy
C0009676|000|hepatic encephalopathy
C0009676|000|septic encephalopathy
C0009676|000|postictal confusion
C0009676|000|icu delirium
C0009676|000|hypoxic encephalopathy
C0009676|000|wernicke’s encephalopathy
C0009676|000|ischemic encephalopathy
C0009676|000|hypoperfusion encephalopathy
C0009676|000|agitated confusion
C0009676|000|restless and confused
C0009676|000|dementia with acute change
C0009676|000|delirium superimposed on dementia
C0009676|000|waxing/waning cognition
C0009676|000|transient confusion
C0009676|000|acute confusional state
C0009676|000|acd (acute confusional disorder)
C0009676|000|delirium nos
C0009676|000|confusional syndrome
C0009676|000|mixed hypoactive/hyperactive delirium
C0009676|000|perplexed
C0009676|000|pocd (postoperative cognitive dysfunction)
C0009676|000|encephalopathic state
C0009676|000|confusional episode
C0009676|000|psycho-organic syndrome
C0009676|000|cognitive impairment
C0009676|000|delirious state
C0009676|000|decreased cognition
C0009676|000|mental confusion
C0009676|000|acute brain dysfunction
C0009676|000|neurocognitive dysfunction
C0009676|000|incoherent
C0009676|000|psychosis (if used for acute confusion)
C0009676|000|muddled
C0009676|000|muddled thinking
C0009676|000|acute brain failure
C0009676|000|disorganized speech
C0009676|000|delayed response
C0009676|000|impaired attention
C0009676|000|short-term memory loss
C0009676|000|unresponsive (when r/t confusion)
C0009676|000|impaired memory and orientation
C0009676|000|reduced arousal
C0009676|000|fluctuating alertness
C0009676|000|depressed level of consciousness
C0009676|000|hyperactive delirium
C0009676|000|hypoactive delirium
C0009676|000|confusional psychosis
C0009676|000|delirium tremens
C0009676|000|delirium due to substance
C0009676|000|withdrawal delirium
C0009676|000|drug-induced confusion
C0009676|000|chemo-induced confusion
C0009676|000|post-stroke confusion
C0009676|000|tia-related confusion
C0009676|000|incoherent mental status
C0009676|000|spoken incoherence
C0009676|000|mistakes place and time
C0009676|000|impaired executive function
C0009676|000|disordered consciousness
C0009676|000|acute brain syndrome
C0009676|000|transient global amnesia (if confused)
C0009676|000|cns dysfunction
C0009676|000|metabolic confusion
C0009676|000|senile confusion
C0009676|000|delirium due to uti
C0009676|000|hospital-acquired delirium
C0009676|000|pod (postoperative delirium)
C0009676|000|encephalopathy nos
C0009676|000|septic confusion
C0009676|000|disorganized behavior
C0009676|000|acute cognitive impairment
C0009676|000|chronic confusion
C0009676|000|substance-induced confusion
C0009676|000|fluctuating cognition
C0009676|000|distractible
C0009676|000|frontal syndrome
C0009676|000|sundowning
C0009676|000|decreased responsiveness
C0009676|000|confusional state nos
C0009676|000|agitated delirium
C0009676|000|restless mental status
C0009676|000|delirium secondary to infection
C0009676|000|delirium of metabolic origin
C0009676|000|delirium due to hypoxia
C0009676|000|paranoia with confusion
C0009676|000|encephalopathic confusion
C0009676|000|mistakes relatives
C0009676|000|word salad
C0009676|000|rambling speech
C0009676|000|unorganized thought process
C0009676|000|thought disorder
C0009676|000|reduced mentation
C0009676|000|abnormal mentation
C0009676|000|periods of unresponsiveness
C0009676|000|clouding of consciousness
C0009676|000|icu psychosis
C0009676|000|acute organic brain syndrome
C0009676|000|toxic psychosis
C0009676|000|organic psychosis
C0009676|000|paranoid confusion
C0009676|000|impaired judgement
C0009676|000|bilious confusion (rare)
C0009676|000|delayed recall
C0009676|000|memory lapses
C0009676|000|impaired cognitive status
C0009676|000|disoriented to time
C0009676|000|disoriented to place
C0009676|000|disoriented to person
C0009676|000|delays in thought
C0009676|000|thought blocking
C0009676|000|forgetful
C0009676|000|attention deficit
C0009676|000|unusual behavior
C0009676|000|disinhibited
C0009676|000|wandering
C0009676|000|not oriented
C0009676|000|not following commands
C0009676|000|memory disturbance
C0009676|000|confabulating
C0009676|000|semantic paraphasia
C0009676|000|aphasic confusion
C0009676|000|acute on chronic confusion
C0009676|000|episodic confusion
C0009676|000|impaired recall
C0009676|000|executive dysfunction
C0009676|000|new cognitive deficit
C0009676|000|fluency disturbance
C0009676|000|paraphasic errors
C0009676|000|confusional arousal
C0009676|000|psychomotor agitation
C0009676|000|psychomotor retardation
C0009676|000|frontal release signs
C0009676|000|amnesia with confusion
C0009676|000|postictal state
C0009676|000|post-ictal confusion
C0009676|000|acute delirium
C0009676|000|dementia with acute confusion
C0009676|000|loc fluctuation
C0009676|000|fluctuating loc
C0009676|000|perseveration (if confused)
C0009676|000|incoherence
C0009676|000|speech disorganization
C0009676|000|language disturbance
C0009676|000|labile mood (if confused)
C0009676|000|inappropriate affect with confusion
C0009676|000|paraphasic confusion
C0009676|000|organically based confusion
C0009676|000|toxic confusion
C0009676|000|leukoencephalopathic confusion
C0009676|000|drug-related encephalopathy
C0009676|000|viral encephalopathy with confusion
C0009676|000|postoperative confusion
C0009676|000|post-anesthesia confusion
C0009676|000|pse (portosystemic encephalopathy)
C0233414|000|impaired attention
C0233414|000|inattentiveness
C0233414|000|poor attention
C0233414|000|decreased attention
C0233414|000|attention deficit
C0233414|000|attention disturbance
C0233414|000|deficit in attention
C0233414|000|distractibility
C0233414|000|difficulty focusing
C0233414|000|shortened attention span
C0233414|000|distraction
C0233414|000|problems concentrating
C0233414|000|concentration deficit
C0233414|000|impaired concentration
C0233414|000|reduced concentration
C0233414|000|decreased concentration
C0233414|000|difficulty concentrating
C0233414|000|unable to concentrate
C0233414|000|concentration disturbance
C0233414|000|attentional impairment
C0233414|000|fluctuating attention
C0233414|000|labile attention
C0233414|000|poor focus
C0233414|000|impaired focus
C0233414|000|easily distracted
C0233414|000|ad
C0233414|000|inability to sustain attention
C0233414|000|inattention
C0233414|000|selective inattention
C0233414|000|failing to attend
C0233414|000|loc impairment (level of consciousness)
C0233414|000|clouded attention
C0233414|000|clouded consciousness
C0233414|000|diffuse attentional disturbance
C0233414|000|nonpersistent attention
C0233414|000|transient attention loss
C0233414|000|brief attention span
C0233414|000|inattentive state
C0233414|000|wandering attention
C0233414|000|unstable attention
C0233414|000|transient inattention
C0233414|000|attention span impairment
C0233414|000|mental inattentiveness
C0233414|000|failure to focus
C0233414|000|short attention span
C0233414|000|distractible
C0233414|000|attentional deficit
C0233414|000|delirium (if used to mean attention disturbance)
C0233414|000|delirious (as shorthand)
C0233414|000|delirium syndrome
C0233414|000|fluctuating awareness
C0233414|000|hypoactive attention
C0233414|000|aao ×3 poor
C0233414|000|impaired vigilance
C0233414|000|reduced vigilance
C0233414|000|dysexecutive syndrome
C0233414|000|executive dysfunction
C0233414|000|non-focal attentional deficit
C0233414|000|subcortical attention impairment
C0233414|000|ischemic attention disturbance
C0233414|000|metabolic attention impairment
C0233414|000|hepatic attention disturbance
C0233414|000|toxic attention impairment
C0233414|000|infectious attention deficit
C0233414|000|delirium d/t infection
C0233414|000|delirium d/t uti
C0233414|000|delirium d/t sepsis
C0233414|000|chemo-induced attention deficit
C0233414|000|attention deficit secondary to tbi
C0233414|000|encephalopathic attention deficit
C0233414|000|drug-induced inattention
C0233414|000|alcohol-related inattention
C0233414|000|paraneoplastic attention deficit
C0233414|000|cancer-related attention deficit
C0233414|000|neurologic attention deficit
C0233414|000|stroke-related inattention
C0233414|000|postictal inattention
C0233414|000|hypoxic attention deficit
C0233414|000|attention deficit – dementia
C0233414|000|vascular attention disturbance
C0233414|000|frontotemporal attention impairment
C0233414|000|alzheimer’s-related inattention
C0233414|000|pd-related inattention
C0233414|000|adhd (in context)
C0233414|000|cognitive slowing
C0233414|000|mental slowing
C0233414|000|bradyphrenia
C0233414|000|psychomotor slowing
C0233414|000|reduced cognitive speed
C0233414|000|attention lapses
C0233414|000|attentional lapses
C0233414|000|fluctuating loc with impaired attention
C0233414|000|impaired divided attention
C0233414|000|poor selective attention
C0233414|000|decreased sustained attention
C0233414|000|impaired sustained attention
C0233414|000|non-sustained attention
C0233414|000|poor task persistence
C0233414|000|vigilance deficit
C0233414|000|monitoring deficit
C0233414|000|reactivity impairment
C0233414|000|impaired responsiveness
C0233414|000|delayed responses
C0233414|000|slow to respond
C0233414|000|diminished alertness
C0233414|000|poor alertness
C0233414|000|reduced mental tracking
C0233414|000|errors in serial 7s
C0233414|000|errors on mmse attention
C0233414|000|failed world backward
C0233414|000|failed serial subtraction
C0233414|000|moca attention deficit
C0233414|000|mmse attention deficit
C0233414|000|consciousness disturbance
C0233414|000|consciousness fluctuation
C0233414|000|encephalopathic state
C0233414|000|encephalopathy with inattention
C0233414|000|cognitive disturbance
C0233414|000|attention-executive dysfunction
C0233414|000|difficulty following conversation
C0233414|000|easily dazed
C0233414|000|mentation fluctuating
C0233414|000|impaired cognitive control
C0233414|000|diffuse cognitive impairment
C0233414|000|loss of vigilance
C0233414|000|decreased mental flexibility
C0233414|000|reduced alertness and attention
C0233414|000|nonverbal inattention
C0233414|000|mild inattentiveness
C0233414|000|moderate inattentiveness
C0233414|000|severe inattentiveness
C0233414|000|attentional failures
C0233414|000|sustained concentration deficit
C0233414|000|task inattention
C0233414|000|slow processing speed
C0233414|000|difficulty maintaining attention
C0233414|000|difficulty with dual tasking
C0233414|000|attention span decreased
C0233414|000|slowed mentation
C0233414|000|impaired mental tracking
C0233414|000|errors on trail making
C0233414|000|omissions on attention tasks
C0233414|000|mental fatigue
C0233414|000|cognitive fatigue
C0233414|000|inattentive subtype
C0233414|000|inattentive presentation
C0454643|000|word finding difficulty
C0454643|000|word-finding difficulty
C0454643|000|word retrieval difficulty
C0454643|000|word finding disorder
C0454643|000|word-finding disorder
C0454643|000|word retrieval deficit
C0454643|000|word-finding deficit
C0454643|000|anomia
C0454643|000|anomic aphasia
C0454643|000|dysnomia
C0454643|000|dysnomia aphasia
C0454643|000|impaired word retrieval
C0454643|000|difficulty with naming
C0454643|000|naming deficit
C0454643|000|naming difficulty
C0454643|000|naming impairment
C0454643|000|impaired naming
C0454643|000|expressive anomia
C0454643|000|aphasia—anomic type
C0454643|000|aphasia (anomic)
C0454643|000|aphasic word-finding difficulty
C0454643|000|aphasic word finding
C0454643|000|aphasic dysnomia
C0454643|000|poststroke anomia
C0454643|000|ischemic anomia
C0454643|000|nonfluent anomia
C0454643|000|fluent anomia
C0454643|000|broca's aphasia with word-finding
C0454643|000|wernicke's aphasia with word-finding
C0454643|000|neurogenic anomia
C0454643|000|vascular anomia
C0454643|000|dementia-related anomia
C0454643|000|ad anomia
C0454643|000|alzheimer's related anomia
C0454643|000|ftd anomia
C0454643|000|semantic anomia
C0454643|000|progressive anomia
C0454643|000|ppa anomia
C0454643|000|primary progressive aphasia with anomia
C0454643|000|tbi-related word-finding
C0454643|000|chemo-induced anomia
C0454643|000|postictal word-finding
C0454643|000|migraine-related word-finding
C0454643|000|tia-related word-finding
C0454643|000|transient anomia
C0454643|000|acute anomia
C0454643|000|chronic anomia
C0454643|000|receptive anomia
C0454643|000|expressive dysnomia
C0454643|000|mild anomic aphasia
C0454643|000|mild word-finding deficit
C0454643|000|moderate word-finding deficit
C0454643|000|severe word-finding impairment
C0454643|000|wfd
C0454643|000|wd
C0454643|000|wfdx
C0454643|000|nfd
C0454643|000|anomic type aphasia
C0454643|000|amnestic aphasia
C0454643|000|loc anomia
C0454643|000|post-op word-finding
C0454643|000|perseverative anomia
C0454643|000|lexical retrieval deficit
C0454643|000|word retrieval impairment
C0454643|000|verbal retrieval deficit
C0454643|000|verbal retrieval impairment
C0454643|000|verbal anomia
C0454643|000|language retrieval deficit
C0454643|000|language retrieval difficulty
C0454643|000|tip-of-the-tongue state
C0454643|000|tot phenomenon
C0454643|000|speech output deficit
C0454643|000|speech hesitation
C0454643|000|lexical-access deficit
C0454643|000|semantic retrieval deficit
C0454643|000|lexical access disorder
C0454643|000|naming latency
C0454643|000|naming hesitation
C0454643|000|naming block
C0454643|000|repetitive anomic errors
C0454643|000|searching for words
C0454643|000|circumlocutory speech
C0454643|000|circumlocution due to anomia
C0454643|000|paraphasic naming errors
C0454643|000|semantic paraphasia (word-finding)
C0454643|000|phonemic paraphasia (word-finding)
C0454643|000|word-finding pauses
C0454643|000|speech arrest (anomia)
C0454643|000|motor aphasia—anomic
C0454643|000|nonfluent aphasia with anomia
C0454643|000|fluent aphasia with anomia
C0454643|000|thalamic anomia
C0454643|000|broca-type word-finding
C0454643|000|wernicke-type word-finding
C0454643|000|global aphasia (with word-finding)
C0454643|000|pca-related anomia
C0454643|000|temporal lobe anomia
C0454643|000|parietal lobe anomia
C0454643|000|frontal lobe anomia
C0454643|000|multifactorial anomia
C0454643|000|amnestic speech
C0454643|000|amnestic disorder with aphasia
C0454643|000|unclassifiable aphasia—anomia dominant
C0454643|000|lbd-related anomia
C0454643|000|vad anomia
C0454643|000|cva anomia
C0454643|000|stroke-related anomia
C0454643|000|sah-related anomia
C0454643|000|functional word-finding
C0454643|000|functional anomia
C0454643|000|psychogenic word-finding issues
C0454643|000|depression-related anomia
C0454643|000|delirium-associated anomia
C0454643|000|delirium word-finding
C0454643|000|focal word-finding deficit
C0454643|000|transient expressive aphasia
C0454643|000|transient expressive anomia
C0454643|000|mild cognitive impairment with anomia
C0454643|000|mci anomia
C0454643|000|age-related word-finding
C0454643|000|developmental anomia
C0454643|000|childhood anomia
C0454643|000|congenital anomia
C0454643|000|genetic anomia
C0454643|000|drug-induced anomia
C0454643|000|medication-induced anomia
C0454643|000|toxic-metabolic word-finding
C0454643|000|metabolic anomia
C0454643|000|encephalopathic anomia
C0454643|000|encephalopathy word-finding
C0454643|000|post-concussive word-finding
C0454643|000|remote word-finding deficit
C0454643|000|hypertensive word-finding
C0454643|000|amyloid anomia
C0454643|000|infectious aphasia—anomic
C0454643|000|autoimmune anomia
C0454643|000|paraneoplastic anomia
C0454643|000|radiation-induced anomia
C0454643|000|postradiation word-finding
C0454643|000|paraphasic speech (anomia)
C0454643|000|mixed aphasia with anomia
C0454643|000|multilingual anomia
C0454643|000|multilingual naming deficit
C0454643|000|secondary anomia
C0454643|000|primary anomia
C0454643|000|acquired anomia
C0454643|000|post-traumatic anomia
C0454643|000|postinfectious word-finding
C0454643|000|postencephalitic anomia
C0454643|000|retograde anomia
C0454643|000|anomic variant ppa
C0454643|000|semantic variant ppa
C0454643|000|logopenic variant ppa with anomia
C0454643|000|logopenic word-finding
C0454643|000|speech disruption (anomic)
C0454643|000|speech disturbance—anomia
C0454643|000|language disturbance—anomia
C0454643|000|pragmatic anomia
C0454643|000|compensated anomia
C0454643|000|residual aphasia—anomic
C0454643|000|remitted aphasia—anomic
C0454643|000|active word-finding deficit
C0454643|000|intermittent word-finding
C0454643|000|cathartic anomia
C0454643|000|verbal access disorder
C0454643|000|lexical semantic deficit
C0454643|000|impaired expressive language (naming)
C0454643|000|aphasia nos (anomic features)
C0454643|000|word-finding issue
C0454643|000|naming problem
C0542476|000|forgetful
C0542476|000|forgetfulness
C0542476|000|memory loss
C0542476|000|memory impairment
C0542476|000|impaired memory
C0542476|000|amnesia
C0542476|000|amnesic
C0542476|000|dementia
C0542476|000|cognitive decline
C0542476|000|cognitive impairment
C0542476|000|dec cognition
C0542476|000|dec memory
C0542476|000|declining memory
C0542476|000|short-term memory loss
C0542476|000|impaired recall
C0542476|000|poor recall
C0542476|000|dec recall
C0542476|000|difficulty remembering
C0542476|000|difficulty recalling
C0542476|000|absent-minded
C0542476|000|absentmindedness
C0542476|000|lapses in memory
C0542476|000|slips of memory
C0542476|000|confused
C0542476|000|confusion
C0542476|000|mental fog
C0542476|000|mentally foggy
C0542476|000|disoriented
C0542476|000|disorientation
C0542476|000|impaired recent memory
C0542476|000|imp rec mem
C0542476|000|impaired remote memory
C0542476|000|imp rem mem
C0542476|000|anterograde amnesia
C0542476|000|retrograde amnesia
C0542476|000|transient global amnesia
C0542476|000|tga
C0542476|000|mnestic deficit
C0542476|000|mnemonic deficit
C0542476|000|forgetting
C0542476|000|trouble remembering
C0542476|000|trouble recalling
C0542476|000|trouble with memory
C0542476|000|stms loss
C0542476|000|ltms loss
C0542476|000|short-term mem loss
C0542476|000|long-term mem loss
C0542476|000|impaired working memory
C0542476|000|deficits in memory
C0542476|000|executive dysfunction
C0542476|000|mild cognitive impairment
C0542476|000|mci
C0542476|000|early dementia
C0542476|000|alzheimer's type memory loss
C0542476|000|ad-type memory loss
C0542476|000|vascular memory impairment
C0542476|000|vascular cognitive impairment
C0542476|000|vci
C0542476|000|post-stroke memory loss
C0542476|000|stroke-related memory loss
C0542476|000|ischemic memory loss
C0542476|000|tbi-related memory loss
C0542476|000|trauma-induced amnesia
C0542476|000|chemobrain
C0542476|000|chemo-induced cognitive impairment
C0542476|000|chemo-induced memory loss
C0542476|000|delirium
C0542476|000|encephalopathic
C0542476|000|encephalopathy-related memory loss
C0542476|000|hiv-associated neurocognitive disorder
C0542476|000|hand
C0542476|000|metabolic memory impairment
C0542476|000|hepatic encephalopathy memory loss
C0542476|000|alcohol-related memory loss
C0542476|000|korsakoff syndrome
C0542476|000|wernicke-korsakoff
C0542476|000|anoxic memory loss
C0542476|000|hypoxic memory loss
C0542476|000|hypoglycemia-related memory loss
C0542476|000|thyroid-related memory impairment
C0542476|000|hypothyroid memory loss
C0542476|000|aging-related memory loss
C0542476|000|age-assoc memory change
C0542476|000|age-assoc mem loss
C0542476|000|senile memory impairment
C0542476|000|senile forgetfulness
C0542476|000|senile dementia
C0542476|000|lewy body-related memory loss
C0542476|000|dlb-associated memory impairment
C0542476|000|frontotemporal memory loss
C0542476|000|ftd-associated memory impairment
C0542476|000|parkinsonian memory impairment
C0542476|000|parkinson's-related memory loss
C0542476|000|pd-associated memory impairment
C0542476|000|ms-related memory impairment
C0542476|000|multiple sclerosis memory loss
C0542476|000|amnestic
C0542476|000|cbi (cognitive behavioral impairment)
C0542476|000|intellectual decline
C0542476|000|progressive memory loss
C0542476|000|transient memory loss
C0542476|000|forgetting names
C0542476|000|forgetting appointments
C0542476|000|repeat questioning
C0542476|000|losing items
C0542476|000|difficulty learning new info
C0542476|000|dysmnestic
C0542476|000|declining cognition
C0542476|000|impaired recognition
C0542476|000|impaired information retention
C0542476|000|impaired learning
C0542476|000|forgetfulness episodes
C0542476|000|episodic memory loss
C0542476|000|impaired autobiographical memory
C0542476|000|poor memory
C0542476|000|dec memory retention
C0542476|000|deficient memory
C0542476|000|suboptimal memory
C0542476|000|slowed mental processing
C0542476|000|impairment in recall
C0542476|000|impaired recent recall
C0542476|000|impaired delayed recall
C0542476|000|inconsistent recall
C0542476|000|diminished memory capacity
C0542476|000|lapses in recall
C0542476|000|poor retention
C0542476|000|memory difficulties
C0542476|000|problems with memory
C0542476|000|diminished short-term memory
C0542476|000|lack of recall
C0542476|000|absent recall
C0542476|000|frontal lobe memory impairment
C0542476|000|temporal lobe memory impairment
C0542476|000|difficulty storing new memories
C0542476|000|working memory difficulty
C0542476|000|amnesia nos
C0542476|000|cognitive deficits
C0542476|000|short term memory impairment
C0542476|000|long term memory impairment
C0542476|000|decline in stm
C0542476|000|decline in ltm
C0542476|000|stm impairment
C0542476|000|ltm impairment
C0542476|000|frequent forgetting
C0542476|000|recurrent memory lapses
C0542476|000|frequent memory lapses
C0542476|000|decreased new learning
C0542476|000|impaired ability to recall facts
C0542476|000|hippocampal memory loss
C0542476|000|executive memory dysfunction
C0542476|000|amnesic episode
C0542476|000|mnestic disturbance
C0542476|000|forgets instructions
C0542476|000|forgetting conversations
C0542476|000|disrupted memory
C0542476|000|amnesic disorder
C0542476|000|amnesic syndrome
C0542476|000|impaired consolidation
C0542476|000|delayed retrieval
C0542476|000|impaired encoding
C0542476|000|imp encoding
C0542476|000|imp retrieval
C0542476|000|impaired retrieval
C1522449|000|radiation therapy
C1522449|000|radiotherapy
C1522449|000|rt
C1522449|000|xrt
C1522449|000|external beam radiation
C1522449|000|external beam rt
C1522449|000|external beam radiotherapy
C1522449|000|ebrt
C1522449|000|radiation tx
C1522449|000|rad tx
C1522449|000|rad therapy
C1522449|000|radio tx
C1522449|000|ionizing radiation therapy
C1522449|000|therapeutic irradiation
C1522449|000|irradiation
C1522449|000|radiotherapeutic procedure
C1522449|000|radiotherapeutics
C1522449|000|radioisotope therapy
C1522449|000|teletherapy
C1522449|000|brachytherapy
C1522449|000|imrt
C1522449|000|intensity-modulated rt
C1522449|000|intensity-modulated radiation therapy
C1522449|000|igrt
C1522449|000|image-guided radiation therapy
C1522449|000|stereotactic radiosurgery
C1522449|000|srs
C1522449|000|sbrt
C1522449|000|stereotactic body radiation therapy
C1522449|000|proton therapy
C1522449|000|proton beam therapy
C1522449|000|pbt
C1522449|000|conventional radiation
C1522449|000|fractionated radiation
C1522449|000|adjuvant rt
C1522449|000|neoadjuvant rt
C1522449|000|conformal rt
C1522449|000|3d crt
C1522449|000|3d conformal radiation
C1522449|000|3d conformal rt
C1522449|000|three-dimensional conformal rt
C1522449|000|pall rt
C1522449|000|palliative radiation
C1522449|000|palliative rt
C1522449|000|whole brain rt
C1522449|000|cns rt
C1522449|000|cranial radiation
C1522449|000|tbi
C1522449|000|total body irradiation
C1522449|000|prophylactic cranial irradiation
C1522449|000|pci
C1522449|000|accelerated rt
C1522449|000|boost radiation
C1522449|000|boost rt
C1522449|000|intraoperative rt
C1522449|000|iort
C1522449|000|rad onc tx
C1522449|000|rad oncology therapy
C1522449|000|radiation course
C1522449|000|external radiation
C1522449|000|radiation
C1522450|000|brachy
C1522451|000|intraop rt
C1522452|000|intraop radiation
C1522453|000|wbrt
C1522454|000|srt
C1522455|000|radiosurgery
C1522456|000|proton
C1522457|000|electron
C1522458|000|photon
C1522459|000|vmat
C1522460|000|volumetric modulated arc radiotherapy
