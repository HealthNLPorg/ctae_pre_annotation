cui|aui|atom_name
C0018801|A0001706|Heart failure
C0018801|A4375418|Heart failure
C0018801|A0418145|HEART FAILURE
C0018801|A9333313|heart failure
C0018801|A4757882|"Heart failure| NOS"
C0018801|A25684844|Failure heart
C0018801|A37223575|Heart Failure
C0018801|A21144613|Cardiac failure
C0018801|A18573120|failure cardiac
C0018801|A9343517|cardiac failure
C0018801|A24668471|Cardiac insufficiency
C0018801|A25735615|Insufficiency cardiac
C0018801|A4394427|cardiac; insufficiency
C0018801|A3319625|Weak heart
C0018801|A0591153|"Weak heart| NOS"
C0018801|A4469213|weak; heart
C0018801|A4419444|heart; insufficiency
C0018801|A22854563|Heart failure NOS (disorder)
C0018801|A32650897|Heart failure
C0018801|A0418147|HEART FAILURE
C0018801|A0418148|HEART FAILURE (NOS)
C0018801|A4386746|heart failure
C0018801|A4782625|Heart failure NOS
C0018801|A1860333|Failure;heart
C0018801|A4413527|failure; heart
C0018801|A23902743|Cardiac Failure
C0018801|A3004656|Cardiac failure
C0018801|A23029834|Weak heart
C0018801|A4765237|"Weak heart| NOS"
C0018801|A18591788|hearts weak
C0018801|A18568810|heart insufficiency
C0018801|A4427526|insufficiency; heart
C0018801|A18647571|heart weakness
C0018801|A1860982|Weakness;heart
C0018801|A22827151|Heart failure (disorder)
C0018801|A4994650|Heart: [weak] or [failure NOS]
C0018801|A23049735|Heart: [weak] or [failure NOS]
C0018801|A0001699|Heart failure
C0018801|A0001703|Heart failure
C0018801|A30071986|Heart failure
C0018801|A32778593|Heart failure
C0018801|A4708533|Heart failure
C0018801|A0411887|FAILURE HEART
C0018801|A22949334|Heart failure NOS
C0018801|A22982915|Heart failure NOS
C0018801|A18573121|failures heart
C0018801|A37232915|Heart Failure
C0018801|A0396685|CARDIAC FAILURE
C0018801|A0540410|"Cardiac failure| NOS"
C0018801|A1257871|Cardiac failure NOS
C0018801|A18698747|insufficiency cardiac
C0018801|A1388938|cardiac insufficiency
C0018801|A8375798|Weak heart
C0018801|A18628924|weak heart
C0018801|A25710455|"Heart failure| unspecified"
C0018801|A1399519|3-16 HEART FAILURE AND OTHER FUNCTIONAL DISORDERS
C0018801|A3488118|Heart failure (disorder)
C0018801|A13947365|cardiac failure (diagnosis)
C0018801|A22953826|Heart: [weak] or [failure NOS] (disorder)
C0018801|A0001704|Heart failure
C0018801|A11973921|Heart failure
C0018801|A30932964|Heart failure
C0018801|A8339687|Heart failure
C0018801|A0714467|Heart failure NOS
C0018801|A16987898|Heart failure NOS
C0018801|A22899326|Heart failure NOS
C0018801|A37225835|Heart Failure
C0018801|A26646995|Cardiac Failure
C0018801|A18610362|cardiac failures
C0018801|A25717599|Cardiac insufficiency
C0018801|A26954697|Cardiac insufficiency
C0018801|A22841831|Insufficiency - cardiac
C0018801|A0568631|"Myocardial failure| NOS"
C0018801|A18554676|myocardial failure
C0018801|A0714471|"Heart failure| unspecified"
C0018801|A0714472|"Heart failure| unspecified"
C0018801|A20107248|"Heart failure| unspecified"
C0018801|A25726900|Heart insufficiency
C0018801|A4419508|heart; weakness
C0018801|A22896578|Heart failure NOS (disorder)
C0018801|A0001701|Heart failure
C0018801|A23873476|Heart failure
C0018801|A25718695|Heart failure
C0018801|A2872568|Heart failure
C0018801|A0480545|heart failure
C0018801|A0556946|"Heart failure| NOS"
C0018801|A8359788|Heart failure NOS
C0018801|A12985263|Heart Failure
C0018801|A4394401|cardiac; failure
C0018801|A4413503|failure; cardiac
C0018801|A18591786|cardiac failure
C0018801|A0396699|CARDIAC INSUFFICIENCY
C0018801|A9334370|cardiac insufficiency
C0018801|A9334797|weak heart
C0018801|A17864489|"Heart failure| unspecified"
C0018801|A1279242|HF - Heart failure
C0018801|A18624576|insufficiency heart
C0018801|A0001700|Heart failure
C0018801|A0001707|Heart failure
C0018801|A17800633|Heart failure
C0018801|A4375419|Heart failure
C0018801|A0418144|HEART FAILURE
C0018801|A21143452|Heart Failure
C0018801|A37374743|Heart Failure
C0018801|A0669023|Cardiac failure
C0018801|A23045758|Cardiac failure NOS
C0018801|A25692337|Cardiac failure NOS
C0018801|A25709267|Cardiac failure (NOS)
C0018801|A1857627|Failure;cardiac
C0018801|A13908563|cardiac failure
C0018801|A0422932|INSUFFICIENCY CARDIAC
C0018801|A0556284|HEART FAILURE AND OTHER FUNCTIONAL DISORDERS
C0018801|A8359789|"Heart failure| unspecified"
C0018801|A25717598|Cardiac function failed
C0018801|A18684586|heart weaknesses
C0018801|A22968943|Heart failure
C0018801|A7191680|Heart failure
C0018801|A0480546|heart failure
C0018801|A18591787|heart failure
C0018801|A18647570|heart failures
C0018801|A2017282|Heart failures
C0018801|A21145427|Cardiac Failure
C0018801|A0396686|CARDIAC FAILURE
C0018801|A4753710|"Cardiac failure| NOS"
C0018801|A8364673|Cardiac failure NOS
C0018801|A23454310|Cardiac insufficiency
C0018801|A18606059|cardiac insufficiency
C0018801|A1857628|Insufficiency;cardiac
C0018801|A22847737|Insufficiency - cardiac
C0018801|A4427487|insufficiency; cardiac
C0018801|A25725745|Cardiac function failure
C0018801|A0480547|heart failure
C0018801|A25685196|Heart failure (NOS)
C0018801|A10782107|Heart Failure
C0018801|A0396687|CARDIAC FAILURE
C0018801|A12032049|Cardiac failure
C0018801|A25692335|Cardiac failure
C0018801|A2849890|Cardiac failure
C0018801|A0396698|CARDIAC INSUFFICIENCY
C0018801|A3280812|HF - Heart failure
